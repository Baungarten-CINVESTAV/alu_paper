// This is the unpowered netlist.
module Top_Module_4_ALU (ALU_Output,
    Exception,
    Operation,
    Overflow,
    Underflow,
    a_operand,
    b_operand);
 output [63:0] ALU_Output;
 output [3:0] Exception;
 input [3:0] Operation;
 output [3:0] Overflow;
 output [3:0] Underflow;
 input [63:0] a_operand;
 input [63:0] b_operand;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05676_ (.I(net12),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05677_ (.I(_01086_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05678_ (.I(_01097_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05679_ (.I(_01108_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05680_ (.I(_01119_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05681_ (.I(_01130_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05682_ (.I(net4),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05683_ (.A1(net3),
    .A2(_01151_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05684_ (.I(net1),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05685_ (.I(net2),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05686_ (.A1(_01173_),
    .A2(_01184_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05687_ (.A1(_01162_),
    .A2(_01195_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05688_ (.I(_01205_),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05689_ (.I(_01216_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05690_ (.I(_01227_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05691_ (.I(_01238_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05692_ (.I(_01130_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05693_ (.I(net76),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05694_ (.I(_01270_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05695_ (.A1(_01260_),
    .A2(_01281_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05696_ (.I(net76),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05697_ (.A1(_01130_),
    .A2(_01303_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05698_ (.I(net2),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05699_ (.A1(net3),
    .A2(_01151_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05700_ (.A1(_01173_),
    .A2(_01336_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05701_ (.A1(_01325_),
    .A2(_01346_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05702_ (.I(_01357_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05703_ (.I(_01368_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05704_ (.I(net1),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05705_ (.I(_01325_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05706_ (.A1(_01390_),
    .A2(_01401_),
    .A3(_01162_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05707_ (.I(_01412_),
    .Z(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05708_ (.I(net3),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05709_ (.I(net4),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05710_ (.I(_01173_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05711_ (.I(_01184_),
    .Z(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05712_ (.A1(_01433_),
    .A2(_01444_),
    .A3(_01455_),
    .A4(_01466_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05713_ (.I(_01477_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05714_ (.A1(_01379_),
    .A2(_01423_),
    .A3(_01488_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05715_ (.A1(_01292_),
    .A2(_01314_),
    .B(_01498_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05716_ (.I(net13),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05717_ (.I(_01520_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05718_ (.I(_01531_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05719_ (.I(_01542_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05720_ (.I(_01553_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05721_ (.I(_01564_),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05722_ (.I(_01575_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05723_ (.I(_01585_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05724_ (.I(net3),
    .ZN(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05725_ (.A1(_01607_),
    .A2(_01444_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05726_ (.A1(_01390_),
    .A2(_01325_),
    .A3(_01618_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05727_ (.I(_01629_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05728_ (.I(_01640_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05729_ (.I(_01651_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05730_ (.A1(_01433_),
    .A2(_01151_),
    .A3(_01455_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05731_ (.A1(_01325_),
    .A2(_01673_),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05732_ (.A1(_01455_),
    .A2(net2),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05733_ (.A1(_01390_),
    .A2(_01184_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05734_ (.A1(_01607_),
    .A2(_01151_),
    .A3(_01694_),
    .A4(_01705_),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05735_ (.A1(_01683_),
    .A2(_01716_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05736_ (.I(_01727_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05737_ (.I(_01281_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05738_ (.I(_01749_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05739_ (.I(_01760_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05740_ (.I(_01770_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05741_ (.I(_01466_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05742_ (.I(_01346_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05743_ (.A1(_01792_),
    .A2(_01803_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05744_ (.I(_01814_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05745_ (.A1(_01433_),
    .A2(_01444_),
    .A3(_01195_),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05746_ (.I(_01836_),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05747_ (.I(_01336_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05748_ (.A1(_01858_),
    .A2(_01705_),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05749_ (.I(_01868_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05750_ (.A1(_01847_),
    .A2(_01879_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05751_ (.A1(_01781_),
    .A2(_01890_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05752_ (.A1(_01825_),
    .A2(_01901_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _05753_ (.A1(_01596_),
    .A2(_01662_),
    .B1(_01738_),
    .B2(_01781_),
    .C1(_01141_),
    .C2(_01912_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05754_ (.A1(_01141_),
    .A2(_01249_),
    .B(_01509_),
    .C(_01923_),
    .ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05755_ (.I(_01401_),
    .Z(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05756_ (.A1(_01433_),
    .A2(_01444_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05757_ (.A1(_01390_),
    .A2(_01944_),
    .A3(_01955_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05758_ (.I(_01966_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05759_ (.I(net77),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05760_ (.I(_01987_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05761_ (.I(_01998_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05762_ (.I(_02009_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05763_ (.A1(_01575_),
    .A2(_02020_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05764_ (.I(_02031_),
    .Z(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05765_ (.I(net29),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05766_ (.I(_02053_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05767_ (.I(net93),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05768_ (.I(_02074_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05769_ (.A1(_02063_),
    .A2(_02085_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05770_ (.I(net26),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05771_ (.I(_02107_),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05772_ (.I(_02118_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05773_ (.I(net90),
    .Z(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05774_ (.I(_02140_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05775_ (.A1(_02129_),
    .A2(_02151_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05776_ (.I(net25),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05777_ (.I(_02172_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05778_ (.I(_02183_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05779_ (.I(_02194_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05780_ (.I(net89),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05781_ (.I(_02216_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05782_ (.I(_02226_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05783_ (.I(_02237_),
    .Z(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05784_ (.A1(_02205_),
    .A2(_02247_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05785_ (.I(net24),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05786_ (.I(_02269_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05787_ (.I(_02280_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05788_ (.I(_02291_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05789_ (.I(net88),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05790_ (.I(_02313_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05791_ (.I(_02324_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05792_ (.A1(_02302_),
    .A2(_02335_),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05793_ (.I(net22),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05794_ (.I(_02357_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05795_ (.I(_02368_),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05796_ (.I(_02379_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05797_ (.I(net86),
    .Z(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05798_ (.I(_02401_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05799_ (.I(_02412_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05800_ (.I(_02423_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05801_ (.A1(_02390_),
    .A2(_02434_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05802_ (.A1(_02390_),
    .A2(_02423_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05803_ (.I(net21),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05804_ (.I(net85),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05805_ (.I(_02478_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05806_ (.I(_02489_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05807_ (.I(_02500_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05808_ (.A1(_02467_),
    .A2(_02510_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05809_ (.I(net20),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05810_ (.I(_02532_),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05811_ (.I(_02543_),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05812_ (.I(_02553_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05813_ (.I(net84),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05814_ (.I(_02575_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05815_ (.I(_02586_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05816_ (.I(_02596_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05817_ (.I(_02607_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05818_ (.A1(_02564_),
    .A2(_02618_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05819_ (.I(net18),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05820_ (.I(_02639_),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05821_ (.I(_02650_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05822_ (.I(_02661_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05823_ (.I(_02672_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05824_ (.I(net82),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05825_ (.I(_02694_),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05826_ (.I(_02704_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05827_ (.I(_02715_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05828_ (.A1(_02683_),
    .A2(_02726_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05829_ (.I(net15),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05830_ (.I(_02748_),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05831_ (.I(_02759_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05832_ (.I(_02769_),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05833_ (.I(_02780_),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05834_ (.I(net79),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05835_ (.I(_02802_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05836_ (.I(_02813_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05837_ (.I(_02824_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05838_ (.I(_02834_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05839_ (.I(_02845_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05840_ (.A1(_02791_),
    .A2(_02856_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05841_ (.I(_02867_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05842_ (.I(net14),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05843_ (.I(_02889_),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05844_ (.I(_02899_),
    .Z(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05845_ (.I(_02910_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05846_ (.I(_02921_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05847_ (.I(net78),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05848_ (.I(_02943_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05849_ (.I(_02954_),
    .Z(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05850_ (.I(_02965_),
    .Z(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05851_ (.I(_02976_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05852_ (.I(_02986_),
    .Z(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05853_ (.A1(_02932_),
    .A2(_02997_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05854_ (.I(_01564_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05855_ (.I(_02020_),
    .Z(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05856_ (.A1(_03019_),
    .A2(_03030_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05857_ (.A1(_01260_),
    .A2(_01281_),
    .B(_02031_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05858_ (.A1(_02932_),
    .A2(_02986_),
    .Z(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05859_ (.A1(_03041_),
    .A2(_03052_),
    .B(_03063_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05860_ (.A1(_02780_),
    .A2(_02834_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05861_ (.A1(_02780_),
    .A2(_02834_),
    .Z(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05862_ (.A1(_03084_),
    .A2(_03095_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05863_ (.A1(_03008_),
    .A2(_03073_),
    .B(_03106_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05864_ (.I(_03030_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05865_ (.A1(_03019_),
    .A2(_03128_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05866_ (.A1(_01292_),
    .A2(_02031_),
    .B(_03139_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05867_ (.A1(_03063_),
    .A2(_03150_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _05868_ (.A1(_02878_),
    .A2(_03117_),
    .B1(_03160_),
    .B2(_03106_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05869_ (.I(net17),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05870_ (.I(_03182_),
    .Z(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05871_ (.I(_03193_),
    .Z(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05872_ (.I(_03204_),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05873_ (.I(_03215_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05874_ (.I(net81),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05875_ (.A1(_03226_),
    .A2(_03237_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05876_ (.I(net81),
    .Z(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05877_ (.I(_03258_),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05878_ (.A1(_03204_),
    .A2(_03269_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05879_ (.A1(_03248_),
    .A2(_03280_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05880_ (.I(_02726_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05881_ (.A1(_02672_),
    .A2(_03302_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05882_ (.I(_03215_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05883_ (.A1(_03324_),
    .A2(_03237_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05884_ (.A1(_03171_),
    .A2(_03291_),
    .B(_03313_),
    .C(_03335_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05885_ (.I(net19),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05886_ (.I(_03356_),
    .Z(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05887_ (.I(_03367_),
    .Z(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05888_ (.I(net83),
    .Z(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05889_ (.I(_03389_),
    .Z(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05890_ (.I(_03400_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05891_ (.A1(_03378_),
    .A2(_03411_),
    .Z(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05892_ (.I(_03356_),
    .Z(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05893_ (.I(net83),
    .Z(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05894_ (.I(_03444_),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05895_ (.A1(_03433_),
    .A2(_03455_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05896_ (.A1(_03422_),
    .A2(_03465_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05897_ (.I(_03378_),
    .Z(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05898_ (.I(_03487_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05899_ (.I(_03411_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05900_ (.A1(_03498_),
    .A2(_03509_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05901_ (.A1(_02737_),
    .A2(_03346_),
    .A3(_03476_),
    .B(_03520_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05902_ (.A1(_02564_),
    .A2(_02618_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05903_ (.I(net21),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05904_ (.I(_03553_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05905_ (.I(_03564_),
    .Z(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05906_ (.I(net85),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05907_ (.A1(_03574_),
    .A2(_03585_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05908_ (.A1(_02629_),
    .A2(_03531_),
    .B(_03542_),
    .C(_03596_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05909_ (.A1(_02456_),
    .A2(_02521_),
    .A3(_03607_),
    .Z(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05910_ (.I(net23),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05911_ (.I(net87),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05912_ (.I(_03640_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05913_ (.I(_03651_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05914_ (.A1(_03629_),
    .A2(_03661_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05915_ (.I(net23),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05916_ (.I(_03683_),
    .Z(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05917_ (.I(_03694_),
    .Z(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05918_ (.I(_03651_),
    .Z(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05919_ (.A1(_03705_),
    .A2(_03716_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05920_ (.A1(_03672_),
    .A2(_03727_),
    .Z(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05921_ (.A1(_03629_),
    .A2(_03716_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05922_ (.A1(_02445_),
    .A2(_03618_),
    .A3(_03738_),
    .B(_03748_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05923_ (.A1(_02302_),
    .A2(_02324_),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05924_ (.I(_03770_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05925_ (.I(_02237_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05926_ (.A1(_02194_),
    .A2(_03792_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05927_ (.A1(_02346_),
    .A2(_03759_),
    .B(_03781_),
    .C(_03803_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05928_ (.I(_02151_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05929_ (.A1(_02129_),
    .A2(_03824_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05930_ (.A1(_02161_),
    .A2(_02258_),
    .A3(_03813_),
    .B(_03835_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05931_ (.I(net28),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05932_ (.I(net92),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05933_ (.I(_03867_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05934_ (.A1(_03856_),
    .A2(_03878_),
    .Z(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05935_ (.I(_03856_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05936_ (.A1(_03900_),
    .A2(_03878_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05937_ (.A1(_03889_),
    .A2(_03911_),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05938_ (.I(_03878_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05939_ (.A1(_03900_),
    .A2(_03933_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05940_ (.A1(_03845_),
    .A2(_03922_),
    .B(_03944_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05941_ (.I(_02063_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05942_ (.A1(_03966_),
    .A2(_02085_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05943_ (.A1(_02096_),
    .A2(_03955_),
    .B(_03977_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05944_ (.I(_03988_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05945_ (.I(_03999_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05946_ (.A1(_01260_),
    .A2(_01781_),
    .B(_03999_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05947_ (.A1(_01314_),
    .A2(_04010_),
    .B(_04021_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05948_ (.A1(_02042_),
    .A2(_04032_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05949_ (.A1(_01976_),
    .A2(_04043_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05950_ (.A1(_01173_),
    .A2(net2),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05951_ (.A1(_01618_),
    .A2(_04065_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05952_ (.I(_04075_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05953_ (.I(_04086_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05954_ (.I(_01749_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05955_ (.A1(_01130_),
    .A2(_04107_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05956_ (.A1(_04118_),
    .A2(_02042_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05957_ (.A1(_04097_),
    .A2(_04129_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05958_ (.I(_01716_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05959_ (.I(_04150_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05960_ (.I(_04161_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05961_ (.A1(_01585_),
    .A2(_03128_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05962_ (.A1(_01858_),
    .A2(_01705_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05963_ (.I(_04193_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05964_ (.I(_04204_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05965_ (.A1(_03128_),
    .A2(_04171_),
    .B1(_04182_),
    .B2(_04215_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05966_ (.A1(_01336_),
    .A2(_04065_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05967_ (.I(_04236_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05968_ (.I(_04247_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05969_ (.I(_04258_),
    .Z(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05970_ (.I(_01216_),
    .Z(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05971_ (.I(_04279_),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05972_ (.I(_02932_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05973_ (.I(_01629_),
    .Z(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05974_ (.I(_04312_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05975_ (.I(_04323_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05976_ (.A1(_04301_),
    .A2(_04334_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05977_ (.A1(_01596_),
    .A2(_04290_),
    .B(_04344_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05978_ (.I(_01673_),
    .Z(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05979_ (.I(_04366_),
    .Z(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05980_ (.I(_04377_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05981_ (.A1(_01792_),
    .A2(_01596_),
    .B(_02042_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05982_ (.A1(_01781_),
    .A2(_01585_),
    .B1(_03128_),
    .B2(_01141_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05983_ (.A1(_04118_),
    .A2(_04182_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05984_ (.A1(_04410_),
    .A2(_04420_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05985_ (.I(_01836_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05986_ (.A1(_04388_),
    .A2(_04399_),
    .B1(_04431_),
    .B2(_04442_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05987_ (.A1(_01141_),
    .A2(_04269_),
    .B(_04355_),
    .C(_04453_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05988_ (.A1(_04054_),
    .A2(_04139_),
    .A3(_04225_),
    .A4(_04464_),
    .ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05989_ (.I(_04086_),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05990_ (.I(_03063_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05991_ (.A1(_04118_),
    .A2(_02042_),
    .B(_04182_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05992_ (.A1(_04495_),
    .A2(_04506_),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05993_ (.A1(_04485_),
    .A2(_04517_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05994_ (.I(_02976_),
    .Z(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05995_ (.A1(_02921_),
    .A2(_04539_),
    .Z(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05996_ (.A1(_04539_),
    .A2(_04171_),
    .B1(_04550_),
    .B2(_04215_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05997_ (.I(_01944_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05998_ (.A1(_04571_),
    .A2(_02997_),
    .B(_04495_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05999_ (.I(_01346_),
    .Z(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06000_ (.I(_04593_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06001_ (.I(_01205_),
    .Z(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06002_ (.I(_04615_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06003_ (.I(_01640_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06004_ (.A1(_02791_),
    .A2(_04637_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06005_ (.A1(_04301_),
    .A2(_04626_),
    .B(_04648_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06006_ (.A1(_01596_),
    .A2(_04269_),
    .B1(_04582_),
    .B2(_04604_),
    .C(_04658_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06007_ (.A1(_03041_),
    .A2(_03052_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06008_ (.I(_03988_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06009_ (.I(_04691_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06010_ (.I(_03988_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06011_ (.A1(_03150_),
    .A2(_04713_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06012_ (.A1(_04680_),
    .A2(_04702_),
    .B(_04724_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06013_ (.A1(_04495_),
    .A2(_04735_),
    .Z(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06014_ (.I(_01477_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06015_ (.A1(_04495_),
    .A2(_04735_),
    .B(_04756_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06016_ (.A1(_01575_),
    .A2(_03030_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06017_ (.A1(_01119_),
    .A2(_04539_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06018_ (.A1(_04778_),
    .A2(_04789_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06019_ (.A1(_01260_),
    .A2(_02997_),
    .A3(_04778_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06020_ (.I(_01270_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06021_ (.A1(_04822_),
    .A2(_02932_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06022_ (.A1(_04800_),
    .A2(_04811_),
    .A3(_04832_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06023_ (.A1(_04800_),
    .A2(_04811_),
    .B(_04832_),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06024_ (.A1(_04420_),
    .A2(_04843_),
    .A3(_04854_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06025_ (.A1(_04843_),
    .A2(_04854_),
    .B(_04420_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06026_ (.A1(_04442_),
    .A2(_04876_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06027_ (.A1(_04745_),
    .A2(_04767_),
    .B1(_04865_),
    .B2(_04887_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06028_ (.A1(_04528_),
    .A2(_04560_),
    .A3(_04669_),
    .A4(_04898_),
    .ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06029_ (.I(_01488_),
    .Z(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06030_ (.I(_04919_),
    .Z(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06031_ (.A1(_03008_),
    .A2(_03073_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06032_ (.I(_03999_),
    .Z(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06033_ (.A1(_04301_),
    .A2(_02997_),
    .B(_03160_),
    .C(_04010_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06034_ (.A1(_04940_),
    .A2(_04951_),
    .B(_04962_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06035_ (.A1(_03106_),
    .A2(_04973_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06036_ (.A1(_02965_),
    .A2(_01564_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06037_ (.A1(_02921_),
    .A2(_02009_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06038_ (.A1(_01119_),
    .A2(_02824_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06039_ (.A1(_04995_),
    .A2(_05006_),
    .A3(_05017_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06040_ (.A1(_01108_),
    .A2(_02976_),
    .A3(_01564_),
    .A4(_02020_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06041_ (.A1(net76),
    .A2(_02769_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06042_ (.A1(_05039_),
    .A2(_05049_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06043_ (.A1(_05028_),
    .A2(_05060_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06044_ (.A1(_04843_),
    .A2(_04865_),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06045_ (.A1(_05071_),
    .A2(_05082_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06046_ (.I(_01847_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06047_ (.I(_05104_),
    .Z(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06048_ (.I(_02954_),
    .Z(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06049_ (.A1(_02910_),
    .A2(_05126_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06050_ (.A1(_03063_),
    .A2(_04506_),
    .B(_05136_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06051_ (.A1(_03106_),
    .A2(_05147_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06052_ (.I(_01216_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06053_ (.I(_05169_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06054_ (.I(_04312_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06055_ (.I(_01401_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06056_ (.I(net15),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06057_ (.I(_05213_),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06058_ (.A1(_05223_),
    .A2(_02813_),
    .Z(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06059_ (.I(_04366_),
    .Z(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06060_ (.A1(_05202_),
    .A2(_05234_),
    .B(_05245_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06061_ (.I(_04247_),
    .Z(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06062_ (.A1(_03324_),
    .A2(_05191_),
    .B1(_03095_),
    .B2(_05256_),
    .C1(_05267_),
    .C2(_04301_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06063_ (.I(_01716_),
    .Z(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06064_ (.I(_05279_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06065_ (.I(_04193_),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06066_ (.I(_05281_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06067_ (.A1(_02845_),
    .A2(_05280_),
    .B1(_05234_),
    .B2(_05282_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06068_ (.A1(_02791_),
    .A2(_05180_),
    .B(_05278_),
    .C(_05283_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06069_ (.A1(_04485_),
    .A2(_05158_),
    .B(_05284_),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06070_ (.A1(_04930_),
    .A2(_04984_),
    .B1(_05093_),
    .B2(_05115_),
    .C(_05285_),
    .ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06071_ (.I(_03291_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06072_ (.I(_05286_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06073_ (.A1(_02878_),
    .A2(_03117_),
    .Z(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06074_ (.I0(_05288_),
    .I1(_03171_),
    .S(_04702_),
    .Z(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06075_ (.A1(_05287_),
    .A2(_05289_),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06076_ (.I(_01966_),
    .Z(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06077_ (.I(_05291_),
    .Z(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06078_ (.A1(_05287_),
    .A2(_05289_),
    .B(_05292_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06079_ (.A1(_01694_),
    .A2(_01955_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06080_ (.I(_05294_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06081_ (.A1(_04865_),
    .A2(_05071_),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06082_ (.A1(_04843_),
    .A2(_05071_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06083_ (.A1(_05028_),
    .A2(_05060_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06084_ (.A1(_05039_),
    .A2(_05049_),
    .B(_05298_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06085_ (.I(_01097_),
    .Z(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06086_ (.A1(_05300_),
    .A2(_03269_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06087_ (.I(_02813_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06088_ (.A1(_05302_),
    .A2(_01542_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06089_ (.A1(_02769_),
    .A2(_02009_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06090_ (.A1(_05136_),
    .A2(_05303_),
    .A3(_05304_),
    .Z(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06091_ (.A1(_05301_),
    .A2(_05305_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06092_ (.A1(_01119_),
    .A2(_02834_),
    .B1(_02976_),
    .B2(_01575_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06093_ (.A1(_04789_),
    .A2(_05303_),
    .B1(_05307_),
    .B2(_05006_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06094_ (.A1(_01270_),
    .A2(_03215_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06095_ (.A1(_05308_),
    .A2(_05309_),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06096_ (.A1(_05306_),
    .A2(_05310_),
    .Z(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06097_ (.A1(_05297_),
    .A2(_05299_),
    .A3(_05311_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06098_ (.A1(_05296_),
    .A2(_05312_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06099_ (.A1(_03095_),
    .A2(_05147_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06100_ (.A1(_03084_),
    .A2(_05314_),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06101_ (.A1(_05287_),
    .A2(_05315_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06102_ (.I(_04086_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06103_ (.I(_02672_),
    .Z(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06104_ (.I(_01683_),
    .Z(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06105_ (.I(_05319_),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06106_ (.I(_01357_),
    .Z(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06107_ (.A1(_03324_),
    .A2(_01227_),
    .B1(_05321_),
    .B2(_05287_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06108_ (.A1(_05318_),
    .A2(_01651_),
    .B1(_03248_),
    .B2(_05320_),
    .C(_05322_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06109_ (.I(_03269_),
    .Z(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06110_ (.I(_05324_),
    .Z(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06111_ (.I(_05279_),
    .Z(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06112_ (.I(net17),
    .Z(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06113_ (.I(net81),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06114_ (.A1(_05327_),
    .A2(_05328_),
    .Z(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06115_ (.I(_05281_),
    .Z(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06116_ (.I(_04236_),
    .Z(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06117_ (.I(_05331_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06118_ (.A1(_05325_),
    .A2(_05326_),
    .B1(_05329_),
    .B2(_05330_),
    .C1(_05332_),
    .C2(_02791_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06119_ (.A1(_05323_),
    .A2(_05333_),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06120_ (.A1(_05295_),
    .A2(_05313_),
    .B1(_05316_),
    .B2(_05317_),
    .C(_05334_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06121_ (.A1(_05290_),
    .A2(_05293_),
    .B(_05335_),
    .ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06122_ (.A1(_02737_),
    .A2(_03313_),
    .Z(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06123_ (.I(_05336_),
    .Z(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06124_ (.A1(_03226_),
    .A2(_05325_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06125_ (.A1(_05288_),
    .A2(_05286_),
    .B(_05338_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06126_ (.A1(_03171_),
    .A2(_05286_),
    .B(_03335_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06127_ (.I0(_05339_),
    .I1(_05340_),
    .S(_04713_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06128_ (.A1(_05337_),
    .A2(_05341_),
    .B(_05291_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06129_ (.A1(_05337_),
    .A2(_05341_),
    .B(_05342_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06130_ (.I(_01847_),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06131_ (.I(_05297_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06132_ (.A1(_05299_),
    .A2(_05311_),
    .Z(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06133_ (.A1(_05299_),
    .A2(_05311_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _06134_ (.A1(_05345_),
    .A2(_05346_),
    .A3(_05347_),
    .B1(_05312_),
    .B2(_04865_),
    .B3(_05071_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06135_ (.A1(_01749_),
    .A2(_03215_),
    .A3(_05308_),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06136_ (.A1(_05306_),
    .A2(_05310_),
    .B(_05349_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06137_ (.A1(_05136_),
    .A2(_05303_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06138_ (.I(_02889_),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06139_ (.I(_05352_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06140_ (.A1(_02813_),
    .A2(_05353_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06141_ (.A1(_05304_),
    .A2(_05351_),
    .B1(_05354_),
    .B2(_04995_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06142_ (.A1(_04822_),
    .A2(_02672_),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06143_ (.A1(_05355_),
    .A2(_05356_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06144_ (.A1(_05301_),
    .A2(_05305_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06145_ (.I(_01086_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06146_ (.I(net82),
    .Z(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06147_ (.A1(_05359_),
    .A2(_05360_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06148_ (.A1(_05324_),
    .A2(_01553_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06149_ (.A1(_05300_),
    .A2(_02715_),
    .A3(_03269_),
    .A4(_01553_),
    .Z(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06150_ (.A1(_05361_),
    .A2(_05362_),
    .B(_05363_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06151_ (.I(_05327_),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06152_ (.A1(_05365_),
    .A2(_01987_),
    .Z(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06153_ (.A1(_02769_),
    .A2(_05126_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06154_ (.A1(_05354_),
    .A2(_05366_),
    .A3(_05367_),
    .Z(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06155_ (.A1(_05364_),
    .A2(_05368_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06156_ (.A1(_05358_),
    .A2(_05369_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06157_ (.A1(_05350_),
    .A2(_05357_),
    .A3(_05370_),
    .Z(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06158_ (.A1(_05346_),
    .A2(_05371_),
    .Z(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06159_ (.A1(_05348_),
    .A2(_05372_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06160_ (.A1(_05348_),
    .A2(_05372_),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06161_ (.I(_04075_),
    .Z(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06162_ (.A1(_03084_),
    .A2(_05314_),
    .B(_05286_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06163_ (.A1(_05329_),
    .A2(_05376_),
    .B(_05336_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06164_ (.A1(_05329_),
    .A2(_05376_),
    .A3(_05337_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06165_ (.A1(_05377_),
    .A2(_05378_),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06166_ (.I(_01868_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06167_ (.A1(_02650_),
    .A2(_02694_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06168_ (.I(_05381_),
    .Z(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06169_ (.A1(_01618_),
    .A2(_01694_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06170_ (.I(_05383_),
    .Z(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06171_ (.A1(_03487_),
    .A2(_04323_),
    .B1(_05384_),
    .B2(_02683_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06172_ (.A1(_05380_),
    .A2(_05382_),
    .B(_05385_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06173_ (.I(_04247_),
    .Z(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06174_ (.A1(_02726_),
    .A2(_04150_),
    .B1(_05387_),
    .B2(_03324_),
    .C1(_05337_),
    .C2(_01803_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06175_ (.A1(_02683_),
    .A2(_01814_),
    .B(_05388_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06176_ (.A1(_05375_),
    .A2(_05379_),
    .B(_05386_),
    .C(_05389_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06177_ (.A1(_05344_),
    .A2(_05373_),
    .A3(_05374_),
    .B(_05390_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06178_ (.A1(_05343_),
    .A2(_05391_),
    .Z(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06179_ (.I(_05392_),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06180_ (.A1(_03422_),
    .A2(_03465_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06181_ (.I(_05393_),
    .Z(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06182_ (.A1(_05318_),
    .A2(_03302_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06183_ (.A1(_03313_),
    .A2(_05339_),
    .B(_05395_),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06184_ (.A1(_02737_),
    .A2(_03346_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06185_ (.I0(_05396_),
    .I1(_05397_),
    .S(_04702_),
    .Z(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06186_ (.A1(_05394_),
    .A2(_05398_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06187_ (.A1(_05394_),
    .A2(_05398_),
    .B(_05292_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06188_ (.A1(_05346_),
    .A2(_05371_),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06189_ (.I(_05401_),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06190_ (.A1(_05402_),
    .A2(_05374_),
    .Z(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06191_ (.A1(_05357_),
    .A2(_05370_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06192_ (.A1(_05350_),
    .A2(_05404_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06193_ (.A1(_05364_),
    .A2(_05368_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06194_ (.I(_02639_),
    .Z(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06195_ (.I(_05407_),
    .Z(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06196_ (.A1(_05408_),
    .A2(_01987_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06197_ (.A1(_03204_),
    .A2(_02954_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06198_ (.A1(_05234_),
    .A2(_05409_),
    .A3(_05410_),
    .Z(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06199_ (.I(_02694_),
    .Z(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06200_ (.I(_01520_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06201_ (.A1(_05412_),
    .A2(_05413_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06202_ (.A1(_03258_),
    .A2(_02899_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06203_ (.A1(_01097_),
    .A2(_03400_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06204_ (.A1(_05414_),
    .A2(_05415_),
    .A3(_05416_),
    .Z(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06205_ (.A1(_05363_),
    .A2(_05411_),
    .A3(_05417_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06206_ (.A1(_05406_),
    .A2(_05418_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06207_ (.A1(_05358_),
    .A2(_05369_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06208_ (.A1(_01270_),
    .A2(_03378_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06209_ (.A1(_05354_),
    .A2(_05367_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06210_ (.A1(_05234_),
    .A2(_04550_),
    .B1(_05366_),
    .B2(_05422_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06211_ (.A1(_05420_),
    .A2(_05421_),
    .A3(_05423_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06212_ (.A1(_04107_),
    .A2(_05318_),
    .A3(_05355_),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06213_ (.A1(_05357_),
    .A2(_05370_),
    .B(_05425_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06214_ (.A1(_05419_),
    .A2(_05424_),
    .A3(_05426_),
    .Z(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06215_ (.A1(_05405_),
    .A2(_05427_),
    .Z(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06216_ (.A1(_05403_),
    .A2(_05428_),
    .Z(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06217_ (.A1(_05394_),
    .A2(_05377_),
    .A3(_05382_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06218_ (.I(_01412_),
    .Z(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06219_ (.A1(_05377_),
    .A2(_05382_),
    .B(_05393_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06220_ (.A1(_05431_),
    .A2(_05432_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06221_ (.I(_02564_),
    .Z(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06222_ (.I(_01640_),
    .Z(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06223_ (.I(_01683_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06224_ (.I(_05436_),
    .Z(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06225_ (.A1(_03487_),
    .A2(_01227_),
    .B1(_05321_),
    .B2(_05394_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06226_ (.A1(_05434_),
    .A2(_05435_),
    .B1(_03422_),
    .B2(_05437_),
    .C(_05438_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06227_ (.A1(_03356_),
    .A2(_03444_),
    .Z(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06228_ (.A1(_03509_),
    .A2(_05326_),
    .B1(_05440_),
    .B2(_05330_),
    .C1(_05332_),
    .C2(_05318_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06229_ (.A1(_05439_),
    .A2(_05441_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06230_ (.A1(_05295_),
    .A2(_05429_),
    .B1(_05430_),
    .B2(_05433_),
    .C(_05442_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06231_ (.A1(_05399_),
    .A2(_05400_),
    .B(_05443_),
    .ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06232_ (.I(_01477_),
    .Z(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06233_ (.I(_05444_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06234_ (.I(_05445_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06235_ (.I(_02564_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06236_ (.A1(_05447_),
    .A2(_02607_),
    .ZN(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06237_ (.A1(_05448_),
    .A2(_03542_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06238_ (.A1(_03498_),
    .A2(_03509_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06239_ (.A1(_05393_),
    .A2(_05396_),
    .B(_05450_),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06240_ (.A1(_04010_),
    .A2(_05451_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06241_ (.A1(_03531_),
    .A2(_04713_),
    .B(_05452_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06242_ (.A1(_05449_),
    .A2(_05453_),
    .ZN(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06243_ (.A1(_05405_),
    .A2(_05427_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06244_ (.I(_05455_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06245_ (.A1(_05402_),
    .A2(_05374_),
    .B(_05428_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06246_ (.A1(_05456_),
    .A2(_05457_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06247_ (.I(_05419_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06248_ (.A1(_05459_),
    .A2(_05424_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06249_ (.A1(_05460_),
    .A2(_05426_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06250_ (.A1(_05459_),
    .A2(_05424_),
    .Z(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06251_ (.A1(_05420_),
    .A2(_05423_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06252_ (.A1(_05420_),
    .A2(_05423_),
    .Z(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06253_ (.A1(_05421_),
    .A2(_05463_),
    .B(_05464_),
    .ZN(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06254_ (.A1(_05300_),
    .A2(_02586_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06255_ (.A1(_05301_),
    .A2(_05414_),
    .Z(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06256_ (.A1(_05467_),
    .A2(_05417_),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06257_ (.A1(_05467_),
    .A2(_05417_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06258_ (.A1(_05411_),
    .A2(_05468_),
    .B(_05469_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06259_ (.A1(_03367_),
    .A2(_01987_),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06260_ (.A1(_03182_),
    .A2(_02802_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06261_ (.A1(_05407_),
    .A2(net78),
    .ZN(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06262_ (.A1(_05472_),
    .A2(_05473_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06263_ (.A1(_05471_),
    .A2(_05474_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06264_ (.A1(net83),
    .A2(net13),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06265_ (.I(_03444_),
    .Z(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06266_ (.A1(_01086_),
    .A2(_05477_),
    .B1(_05360_),
    .B2(_01531_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06267_ (.A1(_05361_),
    .A2(_05476_),
    .B1(_05478_),
    .B2(_05415_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06268_ (.A1(net81),
    .A2(net15),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06269_ (.A1(net82),
    .A2(_05352_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06270_ (.A1(_05476_),
    .A2(_05480_),
    .A3(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06271_ (.A1(_05479_),
    .A2(_05482_),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06272_ (.A1(_05475_),
    .A2(_05483_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06273_ (.I(_05484_),
    .Z(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06274_ (.A1(_05466_),
    .A2(_05470_),
    .A3(_05485_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06275_ (.A1(_04822_),
    .A2(_02553_),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06276_ (.A1(_05406_),
    .A2(_05418_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06277_ (.A1(_03084_),
    .A2(_05410_),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06278_ (.A1(_05409_),
    .A2(_05489_),
    .B1(_05472_),
    .B2(_05367_),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06279_ (.A1(_05488_),
    .A2(_05490_),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06280_ (.A1(_05486_),
    .A2(_05487_),
    .A3(_05491_),
    .Z(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06281_ (.A1(_05462_),
    .A2(_05465_),
    .A3(_05492_),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06282_ (.A1(_05461_),
    .A2(_05493_),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06283_ (.A1(_05458_),
    .A2(_05494_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06284_ (.I(_05104_),
    .Z(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06285_ (.I(_01727_),
    .Z(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06286_ (.I(_05497_),
    .Z(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06287_ (.A1(_05440_),
    .A2(_05432_),
    .A3(_05449_),
    .Z(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06288_ (.A1(_05440_),
    .A2(_05432_),
    .B(_05449_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06289_ (.A1(_05499_),
    .A2(_05500_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06290_ (.I(_04075_),
    .Z(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06291_ (.I(_05502_),
    .Z(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06292_ (.I(_05383_),
    .Z(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06293_ (.I(_05504_),
    .Z(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06294_ (.I(_04247_),
    .Z(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06295_ (.I(_05506_),
    .Z(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06296_ (.A1(_05447_),
    .A2(_05505_),
    .B1(_05507_),
    .B2(_03487_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06297_ (.I(_03574_),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06298_ (.I(_01629_),
    .Z(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06299_ (.I(_05510_),
    .Z(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06300_ (.I(_05281_),
    .Z(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06301_ (.A1(net20),
    .A2(net84),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06302_ (.I(_05513_),
    .Z(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06303_ (.I(_05514_),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06304_ (.A1(_05509_),
    .A2(_05511_),
    .B1(_05512_),
    .B2(_05515_),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06305_ (.I(_05436_),
    .Z(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06306_ (.A1(_01466_),
    .A2(_01673_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06307_ (.I(_05518_),
    .Z(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06308_ (.I(_05519_),
    .Z(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06309_ (.A1(_05434_),
    .A2(_05517_),
    .B1(_05520_),
    .B2(_05449_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06310_ (.A1(_05508_),
    .A2(_05516_),
    .A3(_05521_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06311_ (.A1(_02607_),
    .A2(_05498_),
    .B1(_05501_),
    .B2(_05503_),
    .C(_05522_),
    .ZN(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06312_ (.A1(_05446_),
    .A2(_05454_),
    .B1(_05495_),
    .B2(_05496_),
    .C(_05523_),
    .ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06313_ (.A1(_02467_),
    .A2(_03585_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06314_ (.A1(_05509_),
    .A2(_02510_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06315_ (.A1(_05524_),
    .A2(_05525_),
    .Z(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06316_ (.I(_05526_),
    .Z(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06317_ (.I(_03999_),
    .Z(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06318_ (.A1(_05434_),
    .A2(_02618_),
    .B1(_05393_),
    .B2(_05396_),
    .C(_05450_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06319_ (.A1(_02629_),
    .A2(_03531_),
    .B(_04951_),
    .C(_03542_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06320_ (.A1(_02629_),
    .A2(_05528_),
    .A3(_05529_),
    .B(_05530_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06321_ (.A1(_05527_),
    .A2(_05531_),
    .Z(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06322_ (.A1(_05527_),
    .A2(_05531_),
    .B(_05292_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06323_ (.A1(_05461_),
    .A2(_05493_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06324_ (.A1(_05456_),
    .A2(_05457_),
    .B(_05494_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06325_ (.A1(_05462_),
    .A2(_05492_),
    .Z(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06326_ (.A1(_05462_),
    .A2(_05492_),
    .Z(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06327_ (.A1(_05465_),
    .A2(_05536_),
    .B(_05537_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06328_ (.A1(_05487_),
    .A2(_05491_),
    .Z(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06329_ (.A1(_05486_),
    .A2(_05539_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06330_ (.A1(_05487_),
    .A2(_05491_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06331_ (.A1(_05488_),
    .A2(_05490_),
    .B(_05541_),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06332_ (.I(_05470_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06333_ (.A1(_05543_),
    .A2(_05484_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06334_ (.A1(_05543_),
    .A2(_05485_),
    .Z(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06335_ (.A1(_05466_),
    .A2(_05544_),
    .A3(_05545_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06336_ (.A1(_01303_),
    .A2(_02467_),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06337_ (.A1(_05472_),
    .A2(_05473_),
    .ZN(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06338_ (.A1(_05471_),
    .A2(_05474_),
    .ZN(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06339_ (.A1(_05548_),
    .A2(_05549_),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06340_ (.A1(_05544_),
    .A2(_05547_),
    .A3(_05550_),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06341_ (.A1(_01108_),
    .A2(_02500_),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06342_ (.A1(_02596_),
    .A2(_01585_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06343_ (.A1(_02478_),
    .A2(_05413_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06344_ (.A1(_05466_),
    .A2(_05554_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06345_ (.A1(_05552_),
    .A2(_05553_),
    .B(_05555_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06346_ (.A1(_05479_),
    .A2(_05482_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06347_ (.A1(_05475_),
    .A2(_05483_),
    .B(_05557_),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06348_ (.A1(_02553_),
    .A2(_02009_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06349_ (.I(_03433_),
    .Z(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06350_ (.A1(_05560_),
    .A2(_02661_),
    .A3(_05302_),
    .A4(_02954_),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06351_ (.A1(_02661_),
    .A2(_05302_),
    .B1(_05126_),
    .B2(_03378_),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06352_ (.A1(_05561_),
    .A2(_05562_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06353_ (.A1(_05559_),
    .A2(_05563_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06354_ (.A1(_05477_),
    .A2(_02899_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06355_ (.A1(_02715_),
    .A2(_02921_),
    .B1(_01553_),
    .B2(_03411_),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06356_ (.A1(_05414_),
    .A2(_05565_),
    .B1(_05566_),
    .B2(_05480_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06357_ (.A1(_05360_),
    .A2(_05223_),
    .ZN(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06358_ (.A1(_05329_),
    .A2(_05565_),
    .A3(_05568_),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06359_ (.A1(_05567_),
    .A2(_05569_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06360_ (.A1(_05564_),
    .A2(_05570_),
    .Z(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06361_ (.A1(_05558_),
    .A2(_05571_),
    .Z(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06362_ (.A1(_05556_),
    .A2(_05572_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06363_ (.A1(_05546_),
    .A2(_05551_),
    .A3(_05573_),
    .Z(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06364_ (.A1(_05540_),
    .A2(_05542_),
    .A3(_05574_),
    .ZN(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06365_ (.A1(_05538_),
    .A2(_05575_),
    .Z(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06366_ (.A1(_05534_),
    .A2(_05535_),
    .B(_05576_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06367_ (.A1(_05534_),
    .A2(_05535_),
    .A3(_05576_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06368_ (.A1(_04442_),
    .A2(_05578_),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06369_ (.A1(_05500_),
    .A2(_05514_),
    .A3(_05527_),
    .Z(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06370_ (.A1(_05500_),
    .A2(_05514_),
    .B(_05527_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06371_ (.A1(_05580_),
    .A2(_05581_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06372_ (.I(_05279_),
    .Z(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06373_ (.A1(_03574_),
    .A2(_02510_),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06374_ (.I(_05519_),
    .Z(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06375_ (.I(_01683_),
    .Z(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06376_ (.A1(_02510_),
    .A2(_05583_),
    .B1(_05584_),
    .B2(_05585_),
    .C(_05586_),
    .ZN(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06377_ (.I(_02379_),
    .Z(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06378_ (.I(_05510_),
    .Z(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06379_ (.I(_05331_),
    .Z(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06380_ (.I(_01868_),
    .Z(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06381_ (.A1(_05509_),
    .A2(_04615_),
    .B1(_05591_),
    .B2(_05584_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06382_ (.A1(_05588_),
    .A2(_05589_),
    .B1(_05590_),
    .B2(_05434_),
    .C(_05592_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06383_ (.A1(_05525_),
    .A2(_05587_),
    .B(_05593_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06384_ (.A1(_05577_),
    .A2(_05579_),
    .B1(_05582_),
    .B2(_05317_),
    .C(_05594_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06385_ (.A1(_05532_),
    .A2(_05533_),
    .B(_05595_),
    .ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06386_ (.A1(_05588_),
    .A2(_02434_),
    .Z(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06387_ (.I(_05526_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06388_ (.A1(_02629_),
    .A2(_05597_),
    .A3(_05529_),
    .B(_03596_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06389_ (.A1(_02521_),
    .A2(_03607_),
    .A3(_04010_),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06390_ (.A1(_04713_),
    .A2(_05598_),
    .B(_05599_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06391_ (.A1(_05596_),
    .A2(_05600_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06392_ (.A1(_05486_),
    .A2(_05539_),
    .A3(_05574_),
    .Z(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06393_ (.A1(_05540_),
    .A2(_05574_),
    .Z(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06394_ (.A1(_05542_),
    .A2(_05603_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06395_ (.A1(_05602_),
    .A2(_05604_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06396_ (.A1(_05543_),
    .A2(_05485_),
    .B(_05550_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06397_ (.A1(_05543_),
    .A2(_05485_),
    .A3(_05550_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06398_ (.A1(_05547_),
    .A2(_05606_),
    .B(_05607_),
    .ZN(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06399_ (.I(_05608_),
    .ZN(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06400_ (.A1(_05546_),
    .A2(_05573_),
    .Z(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06401_ (.A1(_05546_),
    .A2(_05573_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06402_ (.A1(_05551_),
    .A2(_05610_),
    .B(_05611_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06403_ (.A1(_05556_),
    .A2(_05572_),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06404_ (.A1(_02575_),
    .A2(_05353_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06405_ (.A1(_01097_),
    .A2(_02412_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06406_ (.A1(_05554_),
    .A2(_05614_),
    .A3(_05615_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06407_ (.A1(_05555_),
    .A2(_05616_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06408_ (.A1(_05567_),
    .A2(_05569_),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06409_ (.A1(_05564_),
    .A2(_05570_),
    .B(_05618_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06410_ (.A1(_05560_),
    .A2(_05302_),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06411_ (.A1(_03564_),
    .A2(_01998_),
    .Z(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06412_ (.A1(_02543_),
    .A2(_05126_),
    .ZN(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06413_ (.A1(_05620_),
    .A2(_05621_),
    .A3(_05622_),
    .ZN(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06414_ (.A1(_03389_),
    .A2(_05223_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06415_ (.A1(_02704_),
    .A2(_02759_),
    .B1(_02910_),
    .B2(_03400_),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06416_ (.A1(_05481_),
    .A2(_05624_),
    .B1(_05625_),
    .B2(_03280_),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06417_ (.A1(_02650_),
    .A2(_05328_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06418_ (.I(_02694_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06419_ (.A1(_05628_),
    .A2(_03193_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06420_ (.A1(_05624_),
    .A2(_05627_),
    .A3(_05629_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06421_ (.A1(_05626_),
    .A2(_05630_),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06422_ (.A1(_05623_),
    .A2(_05631_),
    .Z(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06423_ (.A1(_05617_),
    .A2(_05619_),
    .A3(_05632_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06424_ (.A1(_05558_),
    .A2(_05571_),
    .Z(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06425_ (.A1(_04822_),
    .A2(_02379_),
    .ZN(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06426_ (.A1(_05559_),
    .A2(_05563_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06427_ (.A1(_05561_),
    .A2(_05636_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06428_ (.A1(_05634_),
    .A2(_05635_),
    .A3(_05637_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06429_ (.A1(_05613_),
    .A2(_05633_),
    .A3(_05638_),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06430_ (.A1(_05609_),
    .A2(_05612_),
    .A3(_05639_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06431_ (.A1(_05538_),
    .A2(_05575_),
    .Z(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06432_ (.A1(_05641_),
    .A2(_05577_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06433_ (.A1(_05605_),
    .A2(_05640_),
    .A3(_05642_),
    .Z(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06434_ (.I(_01727_),
    .Z(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06435_ (.A1(_05524_),
    .A2(_05581_),
    .A3(_05596_),
    .Z(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06436_ (.A1(_05524_),
    .A2(_05581_),
    .B(_05596_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06437_ (.A1(_05645_),
    .A2(_05646_),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06438_ (.I(_05502_),
    .Z(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06439_ (.A1(_02390_),
    .A2(_05505_),
    .B1(_05507_),
    .B2(_05509_),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06440_ (.I(_03705_),
    .Z(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06441_ (.A1(_02379_),
    .A2(_02434_),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06442_ (.I(_05651_),
    .Z(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06443_ (.I(_05652_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06444_ (.A1(_05650_),
    .A2(_05511_),
    .B1(_05512_),
    .B2(_05653_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06445_ (.A1(_05588_),
    .A2(_05517_),
    .B1(_05520_),
    .B2(_05596_),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06446_ (.A1(_05649_),
    .A2(_05654_),
    .A3(_05655_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06447_ (.A1(_02434_),
    .A2(_05644_),
    .B1(_05647_),
    .B2(_05648_),
    .C(_05656_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06448_ (.A1(_05446_),
    .A2(_05601_),
    .B1(_05643_),
    .B2(_05496_),
    .C(_05657_),
    .ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06449_ (.A1(_02445_),
    .A2(_03618_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06450_ (.A1(_02456_),
    .A2(_05598_),
    .B(_02445_),
    .ZN(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06451_ (.A1(_04702_),
    .A2(_05659_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06452_ (.A1(_05658_),
    .A2(_05528_),
    .B(_05660_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06453_ (.A1(_03738_),
    .A2(_05661_),
    .Z(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06454_ (.I(_05291_),
    .Z(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06455_ (.A1(_03738_),
    .A2(_05661_),
    .B(_05663_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06456_ (.I(_05294_),
    .Z(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06457_ (.I(_05665_),
    .Z(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06458_ (.A1(_05612_),
    .A2(_05639_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06459_ (.A1(_05612_),
    .A2(_05639_),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06460_ (.A1(_05609_),
    .A2(_05667_),
    .B(_05668_),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06461_ (.A1(_05561_),
    .A2(_05636_),
    .A3(_05634_),
    .ZN(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06462_ (.A1(_05561_),
    .A2(_05636_),
    .B(_05634_),
    .ZN(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06463_ (.A1(_05635_),
    .A2(_05670_),
    .B(_05671_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06464_ (.A1(_05556_),
    .A2(_05572_),
    .B(_05633_),
    .ZN(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06465_ (.A1(_05556_),
    .A2(_05572_),
    .A3(_05633_),
    .ZN(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06466_ (.A1(_05673_),
    .A2(_05638_),
    .B(_05674_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06467_ (.A1(_05619_),
    .A2(_05632_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06468_ (.A1(_05617_),
    .A2(_00000_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06469_ (.A1(_01086_),
    .A2(_03640_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06470_ (.A1(_02412_),
    .A2(_05413_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06471_ (.A1(_05300_),
    .A2(_02423_),
    .B1(_02500_),
    .B2(_01542_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06472_ (.A1(_05552_),
    .A2(_00003_),
    .B1(_00004_),
    .B2(_05614_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06473_ (.A1(_02575_),
    .A2(_02759_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06474_ (.A1(_02489_),
    .A2(_02910_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06475_ (.A1(_00003_),
    .A2(_00006_),
    .A3(_00007_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06476_ (.A1(_00005_),
    .A2(_00008_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06477_ (.A1(_00002_),
    .A2(_00009_),
    .Z(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06478_ (.A1(_05626_),
    .A2(_05630_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06479_ (.A1(_05623_),
    .A2(_05631_),
    .B(_00011_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06480_ (.A1(_05555_),
    .A2(_05616_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06481_ (.A1(net20),
    .A2(net79),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06482_ (.A1(net22),
    .A2(net77),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06483_ (.A1(net21),
    .A2(_02943_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06484_ (.A1(_00014_),
    .A2(_00015_),
    .A3(_00016_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06485_ (.A1(_03444_),
    .A2(_03182_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06486_ (.A1(_05360_),
    .A2(_03193_),
    .B1(_05223_),
    .B2(_05477_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06487_ (.A1(_05568_),
    .A2(_00018_),
    .B1(_00019_),
    .B2(_05627_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06488_ (.A1(_03433_),
    .A2(_03258_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06489_ (.A1(_05381_),
    .A2(_00018_),
    .A3(_00021_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06490_ (.A1(_00017_),
    .A2(_00020_),
    .A3(_00022_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06491_ (.A1(_00013_),
    .A2(_00023_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06492_ (.A1(_00012_),
    .A2(_00024_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06493_ (.A1(_00010_),
    .A2(_00025_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06494_ (.A1(_05619_),
    .A2(_05632_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06495_ (.A1(_01281_),
    .A2(_03705_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06496_ (.A1(_05620_),
    .A2(_05622_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06497_ (.A1(_05620_),
    .A2(_05622_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06498_ (.A1(_05621_),
    .A2(_00029_),
    .B(_00030_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06499_ (.A1(_00027_),
    .A2(_00028_),
    .A3(_00031_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06500_ (.A1(_00001_),
    .A2(_00026_),
    .A3(_00032_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06501_ (.A1(_05675_),
    .A2(_00033_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06502_ (.A1(_05672_),
    .A2(_00034_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06503_ (.A1(_05669_),
    .A2(_00035_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06504_ (.I(_05640_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06505_ (.A1(_05605_),
    .A2(_00037_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06506_ (.A1(_05641_),
    .A2(_05577_),
    .B1(_05605_),
    .B2(_00037_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06507_ (.A1(_00038_),
    .A2(_00039_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06508_ (.I(_00040_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06509_ (.A1(_00036_),
    .A2(_00041_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06510_ (.A1(_03672_),
    .A2(_03727_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06511_ (.A1(_00043_),
    .A2(_05646_),
    .A3(_05652_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06512_ (.I(_01412_),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06513_ (.A1(_05646_),
    .A2(_05652_),
    .B(_00043_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06514_ (.A1(_00045_),
    .A2(_00046_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06515_ (.I(_02291_),
    .Z(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06516_ (.I(_01216_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06517_ (.A1(_05650_),
    .A2(_00049_),
    .B1(_01368_),
    .B2(_00043_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06518_ (.A1(_00048_),
    .A2(_05435_),
    .B1(_03672_),
    .B2(_05437_),
    .C(_00050_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06519_ (.A1(_03629_),
    .A2(_03661_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06520_ (.A1(_03716_),
    .A2(_05326_),
    .B1(_00052_),
    .B2(_05330_),
    .C1(_05332_),
    .C2(_05588_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06521_ (.A1(_00051_),
    .A2(_00053_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06522_ (.A1(_05666_),
    .A2(_00042_),
    .B1(_00044_),
    .B2(_00047_),
    .C(_00054_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06523_ (.A1(_05662_),
    .A2(_05664_),
    .B(_00055_),
    .ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06524_ (.A1(_02346_),
    .A2(_03770_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06525_ (.A1(_05650_),
    .A2(_03661_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06526_ (.A1(_03738_),
    .A2(_05659_),
    .B(_00057_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06527_ (.I0(_00058_),
    .I1(_03759_),
    .S(_04691_),
    .Z(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06528_ (.A1(_00056_),
    .A2(_00059_),
    .Z(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06529_ (.A1(_05669_),
    .A2(_00035_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06530_ (.A1(_00036_),
    .A2(_00041_),
    .B(_00061_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06531_ (.A1(_05675_),
    .A2(_00033_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06532_ (.A1(_05672_),
    .A2(_00034_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06533_ (.A1(_00063_),
    .A2(_00064_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06534_ (.A1(_00027_),
    .A2(_00031_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06535_ (.A1(_00027_),
    .A2(_00031_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06536_ (.A1(_00028_),
    .A2(_00066_),
    .B(_00067_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06537_ (.A1(_00001_),
    .A2(_00026_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06538_ (.A1(_00028_),
    .A2(_00066_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06539_ (.A1(_00001_),
    .A2(_00026_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06540_ (.A1(_00069_),
    .A2(_00070_),
    .B(_00071_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06541_ (.A1(_01760_),
    .A2(_02280_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06542_ (.A1(_00013_),
    .A2(_00023_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06543_ (.A1(_00012_),
    .A2(_00024_),
    .B(_00074_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06544_ (.A1(_00014_),
    .A2(_00016_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06545_ (.A1(net21),
    .A2(net79),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06546_ (.A1(_05622_),
    .A2(_00077_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06547_ (.A1(_00015_),
    .A2(_00076_),
    .B(_00078_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06548_ (.A1(_00075_),
    .A2(_00079_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06549_ (.A1(_00073_),
    .A2(_00080_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06550_ (.A1(_00010_),
    .A2(_00025_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06551_ (.A1(_00002_),
    .A2(_00009_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06552_ (.A1(_00020_),
    .A2(_00022_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06553_ (.A1(_00020_),
    .A2(_00022_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06554_ (.A1(_00017_),
    .A2(_00084_),
    .B(_00085_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06555_ (.A1(_00005_),
    .A2(_00008_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06556_ (.A1(net23),
    .A2(net77),
    .Z(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06557_ (.A1(_02357_),
    .A2(_02943_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06558_ (.A1(_00077_),
    .A2(_00088_),
    .A3(_00089_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06559_ (.A1(_05408_),
    .A2(_05628_),
    .B1(_03193_),
    .B2(_05477_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06560_ (.A1(_03389_),
    .A2(_05407_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06561_ (.A1(_00021_),
    .A2(_00091_),
    .B1(_00092_),
    .B2(_05629_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06562_ (.A1(_02532_),
    .A2(_05328_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06563_ (.A1(_03433_),
    .A2(_05412_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06564_ (.A1(_00092_),
    .A2(_00094_),
    .A3(_00095_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06565_ (.A1(_00090_),
    .A2(_00093_),
    .A3(_00096_),
    .Z(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06566_ (.A1(_00087_),
    .A2(_00097_),
    .Z(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06567_ (.A1(_00086_),
    .A2(_00098_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06568_ (.A1(_05359_),
    .A2(_02313_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06569_ (.A1(_03661_),
    .A2(_03019_),
    .B(_00100_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06570_ (.A1(_02313_),
    .A2(_01531_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06571_ (.A1(_00002_),
    .A2(_00102_),
    .Z(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06572_ (.I(_00103_),
    .Z(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06573_ (.A1(_00101_),
    .A2(_00104_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06574_ (.A1(_02412_),
    .A2(_05353_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06575_ (.A1(_00003_),
    .A2(_00007_),
    .Z(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06576_ (.A1(_05554_),
    .A2(_00106_),
    .B1(_00107_),
    .B2(_00006_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06577_ (.A1(_02586_),
    .A2(_05365_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06578_ (.A1(_02489_),
    .A2(_02759_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06579_ (.A1(_00106_),
    .A2(_00109_),
    .A3(_00110_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06580_ (.A1(_00108_),
    .A2(_00111_),
    .Z(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06581_ (.A1(_00105_),
    .A2(_00112_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06582_ (.A1(_00083_),
    .A2(_00099_),
    .A3(_00113_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06583_ (.A1(_00082_),
    .A2(_00114_),
    .Z(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06584_ (.A1(_00081_),
    .A2(_00115_),
    .Z(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06585_ (.A1(_00068_),
    .A2(_00072_),
    .A3(_00116_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06586_ (.I(_00117_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06587_ (.A1(_00065_),
    .A2(_00118_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06588_ (.A1(_00063_),
    .A2(_00064_),
    .A3(_00117_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06589_ (.A1(_00119_),
    .A2(_00120_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06590_ (.A1(_00062_),
    .A2(_00121_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06591_ (.A1(_00052_),
    .A2(_00046_),
    .A3(_00056_),
    .Z(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06592_ (.A1(_00052_),
    .A2(_00046_),
    .B(_00056_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06593_ (.A1(_00123_),
    .A2(_00124_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06594_ (.I(_05387_),
    .Z(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06595_ (.A1(_05650_),
    .A2(_00126_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06596_ (.A1(_00048_),
    .A2(_02335_),
    .A3(_05282_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06597_ (.I(_02194_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06598_ (.I(_05510_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06599_ (.I(_05504_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06600_ (.A1(_00129_),
    .A2(_00130_),
    .B1(_00131_),
    .B2(_02302_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06601_ (.I(_05518_),
    .Z(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06602_ (.A1(_00048_),
    .A2(_05319_),
    .B1(_00133_),
    .B2(_00056_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06603_ (.A1(_00127_),
    .A2(_00128_),
    .A3(_00132_),
    .A4(_00134_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06604_ (.A1(_02335_),
    .A2(_05644_),
    .B1(_00125_),
    .B2(_05648_),
    .C(_00135_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06605_ (.A1(_05446_),
    .A2(_00060_),
    .B1(_00122_),
    .B2(_05496_),
    .C(_00136_),
    .ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06606_ (.I(_01488_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06607_ (.I(_00137_),
    .Z(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06608_ (.A1(_02205_),
    .A2(_02247_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06609_ (.I(_00139_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06610_ (.I(_02346_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06611_ (.A1(_03770_),
    .A2(_00058_),
    .B(_00141_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06612_ (.A1(_00140_),
    .A2(_00142_),
    .Z(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06613_ (.A1(_02346_),
    .A2(_03759_),
    .B(_03781_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06614_ (.A1(_00144_),
    .A2(_00140_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06615_ (.I0(_00143_),
    .I1(_00145_),
    .S(_05528_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06616_ (.A1(_00036_),
    .A2(_00119_),
    .A3(_00120_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06617_ (.A1(_00061_),
    .A2(_00120_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06618_ (.A1(_00040_),
    .A2(_00147_),
    .B(_00148_),
    .C(_00119_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06619_ (.A1(_00072_),
    .A2(_00116_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06620_ (.A1(_00072_),
    .A2(_00116_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06621_ (.A1(_00068_),
    .A2(_00150_),
    .B(_00151_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06622_ (.A1(_01770_),
    .A2(_02291_),
    .A3(_00080_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06623_ (.A1(_00075_),
    .A2(_00079_),
    .B(_00153_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06624_ (.A1(_00010_),
    .A2(_00025_),
    .A3(_00114_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06625_ (.A1(_00081_),
    .A2(_00115_),
    .B(_00155_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06626_ (.A1(_04107_),
    .A2(_02183_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06627_ (.A1(_00087_),
    .A2(_00097_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06628_ (.A1(_00086_),
    .A2(_00098_),
    .B(_00158_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06629_ (.A1(_00077_),
    .A2(_00089_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06630_ (.A1(net22),
    .A2(net79),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06631_ (.A1(_00016_),
    .A2(_00161_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06632_ (.A1(_00088_),
    .A2(_00160_),
    .B(_00162_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06633_ (.A1(_00159_),
    .A2(_00163_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06634_ (.A1(_00157_),
    .A2(_00164_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06635_ (.A1(_00083_),
    .A2(_00113_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06636_ (.A1(_00083_),
    .A2(_00113_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06637_ (.A1(_00099_),
    .A2(_00166_),
    .B(_00167_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06638_ (.A1(_00101_),
    .A2(_00104_),
    .A3(_00112_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06639_ (.A1(_03640_),
    .A2(_05353_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06640_ (.A1(_01108_),
    .A2(_02237_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06641_ (.A1(_00102_),
    .A2(_00170_),
    .A3(_00171_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06642_ (.A1(net86),
    .A2(_05213_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06643_ (.A1(_00106_),
    .A2(_00110_),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06644_ (.A1(_00007_),
    .A2(_00173_),
    .B1(_00174_),
    .B2(_00109_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06645_ (.A1(net84),
    .A2(net18),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06646_ (.A1(net85),
    .A2(_03182_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06647_ (.A1(_00173_),
    .A2(_00176_),
    .A3(_00177_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06648_ (.A1(_00103_),
    .A2(_00178_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06649_ (.A1(_00175_),
    .A2(_00179_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06650_ (.A1(_00172_),
    .A2(_00180_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06651_ (.A1(_00169_),
    .A2(_00181_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06652_ (.A1(_00093_),
    .A2(_00096_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06653_ (.A1(_00093_),
    .A2(_00096_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06654_ (.A1(_00090_),
    .A2(_00183_),
    .B(_00184_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06655_ (.A1(_00108_),
    .A2(_00111_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06656_ (.A1(net24),
    .A2(net77),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06657_ (.A1(_03683_),
    .A2(net78),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06658_ (.A1(_00161_),
    .A2(_00187_),
    .A3(_00188_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06659_ (.I(_00189_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06660_ (.A1(_03455_),
    .A2(_05408_),
    .B1(_05412_),
    .B2(_03367_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06661_ (.A1(_03465_),
    .A2(_05382_),
    .B1(_00094_),
    .B2(_00191_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06662_ (.A1(_03553_),
    .A2(_05328_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06663_ (.A1(_02532_),
    .A2(_05412_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06664_ (.A1(_05440_),
    .A2(_00193_),
    .A3(_00194_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06665_ (.A1(_00190_),
    .A2(_00192_),
    .A3(_00195_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06666_ (.A1(_00186_),
    .A2(_00196_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06667_ (.A1(_00185_),
    .A2(_00197_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06668_ (.A1(_00182_),
    .A2(_00198_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06669_ (.A1(_00168_),
    .A2(_00199_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06670_ (.A1(_00165_),
    .A2(_00200_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06671_ (.A1(_00156_),
    .A2(_00201_),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06672_ (.A1(_00154_),
    .A2(_00202_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06673_ (.A1(_00152_),
    .A2(_00203_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06674_ (.A1(_00149_),
    .A2(_00204_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06675_ (.A1(_02291_),
    .A2(_02335_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06676_ (.A1(_00140_),
    .A2(_00124_),
    .A3(_00206_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06677_ (.A1(_00124_),
    .A2(_00206_),
    .B(_00139_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06678_ (.A1(_00207_),
    .A2(_00208_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06679_ (.I(_02118_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06680_ (.I(_04312_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06681_ (.I(_05331_),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06682_ (.I(_01466_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06683_ (.A1(_00213_),
    .A2(_02247_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06684_ (.A1(_00140_),
    .A2(_00214_),
    .B(_05245_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06685_ (.A1(_00210_),
    .A2(_00211_),
    .B1(_00212_),
    .B2(_00048_),
    .C(_00215_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06686_ (.I(_05279_),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06687_ (.A1(_02205_),
    .A2(_03792_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06688_ (.A1(_02247_),
    .A2(_00217_),
    .B1(_00218_),
    .B2(_05330_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06689_ (.A1(_00129_),
    .A2(_04290_),
    .B(_00216_),
    .C(_00219_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06690_ (.A1(_05666_),
    .A2(_00205_),
    .B1(_00209_),
    .B2(_05317_),
    .C(_00220_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06691_ (.A1(_00138_),
    .A2(_00146_),
    .B(_00221_),
    .ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06692_ (.A1(_02118_),
    .A2(_03824_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06693_ (.A1(_00129_),
    .A2(_03792_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06694_ (.A1(_00223_),
    .A2(_00142_),
    .B(_03803_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06695_ (.A1(_02258_),
    .A2(_03813_),
    .B(_04691_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06696_ (.A1(_04951_),
    .A2(_00224_),
    .B(_00225_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06697_ (.A1(_00222_),
    .A2(_00226_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06698_ (.A1(_00218_),
    .A2(_00208_),
    .A3(_00222_),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06699_ (.A1(_00218_),
    .A2(_00208_),
    .B(_00222_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06700_ (.A1(_05375_),
    .A2(_00228_),
    .A3(_00229_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06701_ (.I(_03900_),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06702_ (.I(_04312_),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06703_ (.I(_00232_),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06704_ (.I(_05384_),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06705_ (.I(_04258_),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06706_ (.A1(_00231_),
    .A2(_00233_),
    .B1(_00234_),
    .B2(_02129_),
    .C1(_00235_),
    .C2(_00129_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06707_ (.I(_05319_),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06708_ (.I(_01803_),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06709_ (.A1(_00210_),
    .A2(_03824_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06710_ (.I(_01716_),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06711_ (.A1(_03824_),
    .A2(_00240_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06712_ (.A1(_05380_),
    .A2(_00239_),
    .B(_00241_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06713_ (.A1(_00210_),
    .A2(_00237_),
    .B1(_00222_),
    .B2(_00238_),
    .C(_00242_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06714_ (.I(_05294_),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06715_ (.A1(_00152_),
    .A2(_00203_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06716_ (.A1(_00149_),
    .A2(_00204_),
    .B(_00245_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06717_ (.A1(_00156_),
    .A2(_00201_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06718_ (.A1(_00154_),
    .A2(_00202_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06719_ (.A1(_01770_),
    .A2(_02194_),
    .A3(_00164_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06720_ (.A1(_00159_),
    .A2(_00163_),
    .B(_00249_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06721_ (.A1(_00168_),
    .A2(_00199_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06722_ (.A1(_00165_),
    .A2(_00200_),
    .B(_00251_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06723_ (.A1(_04107_),
    .A2(_02107_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06724_ (.A1(_00186_),
    .A2(_00196_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06725_ (.A1(_00185_),
    .A2(_00197_),
    .B(_00254_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06726_ (.A1(_00161_),
    .A2(_00188_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06727_ (.A1(_03683_),
    .A2(_02802_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06728_ (.A1(_00089_),
    .A2(_00257_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06729_ (.A1(_00187_),
    .A2(_00256_),
    .B(_00258_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06730_ (.A1(_00255_),
    .A2(_00259_),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06731_ (.A1(_00253_),
    .A2(_00260_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06732_ (.A1(_00101_),
    .A2(_00104_),
    .A3(_00112_),
    .A4(_00181_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06733_ (.A1(_00182_),
    .A2(_00198_),
    .B(_00262_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06734_ (.A1(_00172_),
    .A2(_00180_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06735_ (.A1(net12),
    .A2(_02140_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06736_ (.A1(net89),
    .A2(_01520_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06737_ (.A1(net87),
    .A2(_05213_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06738_ (.I(net88),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06739_ (.A1(_00268_),
    .A2(_05352_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06740_ (.A1(_00266_),
    .A2(_00267_),
    .A3(_00269_),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06741_ (.A1(_00265_),
    .A2(_00270_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06742_ (.A1(_00173_),
    .A2(_00177_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06743_ (.A1(_02401_),
    .A2(net17),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06744_ (.A1(_00110_),
    .A2(_00273_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06745_ (.A1(_00176_),
    .A2(_00272_),
    .B(_00274_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06746_ (.A1(_05359_),
    .A2(_02226_),
    .B1(_02313_),
    .B2(_01542_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06747_ (.A1(_00100_),
    .A2(_00266_),
    .B1(_00276_),
    .B2(_00170_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06748_ (.A1(net84),
    .A2(net19),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06749_ (.A1(_02478_),
    .A2(_02650_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06750_ (.A1(_00273_),
    .A2(_00278_),
    .A3(_00279_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06751_ (.A1(_00277_),
    .A2(_00280_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06752_ (.A1(_00275_),
    .A2(_00281_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06753_ (.A1(_00271_),
    .A2(_00282_),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06754_ (.A1(_00192_),
    .A2(_00195_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06755_ (.A1(_00192_),
    .A2(_00195_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06756_ (.A1(_00190_),
    .A2(_00284_),
    .B(_00285_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06757_ (.A1(_00104_),
    .A2(_00178_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06758_ (.A1(_00103_),
    .A2(_00178_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06759_ (.A1(_00175_),
    .A2(_00287_),
    .B(_00288_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06760_ (.A1(_02172_),
    .A2(_01998_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06761_ (.A1(net24),
    .A2(net78),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06762_ (.A1(_00257_),
    .A2(_00291_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06763_ (.A1(_00290_),
    .A2(_00292_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06764_ (.A1(_03465_),
    .A2(_00194_),
    .Z(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06765_ (.A1(_02543_),
    .A2(_03455_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06766_ (.A1(_00193_),
    .A2(_00294_),
    .B1(_00295_),
    .B2(_00095_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06767_ (.A1(_02368_),
    .A2(_03258_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06768_ (.A1(_03564_),
    .A2(_02704_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06769_ (.A1(_00295_),
    .A2(_00297_),
    .A3(_00298_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06770_ (.A1(_00293_),
    .A2(_00296_),
    .A3(_00299_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06771_ (.A1(_00286_),
    .A2(_00289_),
    .A3(_00300_),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06772_ (.A1(_00264_),
    .A2(_00283_),
    .A3(_00301_),
    .Z(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06773_ (.A1(_00263_),
    .A2(_00302_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06774_ (.A1(_00261_),
    .A2(_00303_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06775_ (.A1(_00252_),
    .A2(_00304_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06776_ (.A1(_00250_),
    .A2(_00305_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06777_ (.A1(_00247_),
    .A2(_00248_),
    .B(_00306_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06778_ (.A1(_00247_),
    .A2(_00248_),
    .A3(_00306_),
    .Z(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06779_ (.A1(_00307_),
    .A2(_00308_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06780_ (.A1(_00246_),
    .A2(_00309_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06781_ (.A1(_00244_),
    .A2(_00310_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06782_ (.A1(_00230_),
    .A2(_00236_),
    .A3(_00243_),
    .A4(_00311_),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06783_ (.A1(_00138_),
    .A2(_00227_),
    .B(_00312_),
    .ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06784_ (.A1(_03835_),
    .A2(_00224_),
    .B(_02161_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06785_ (.A1(_04691_),
    .A2(_00313_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06786_ (.A1(_03845_),
    .A2(_04951_),
    .B(_00314_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06787_ (.A1(_03922_),
    .A2(_00315_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06788_ (.A1(_00149_),
    .A2(_00204_),
    .A3(_00309_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06789_ (.A1(_00247_),
    .A2(_00248_),
    .A3(_00306_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06790_ (.A1(_00245_),
    .A2(_00307_),
    .B(_00318_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06791_ (.A1(_00317_),
    .A2(_00319_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06792_ (.A1(_00252_),
    .A2(_00304_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06793_ (.A1(_00250_),
    .A2(_00305_),
    .B(_00321_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06794_ (.A1(_01770_),
    .A2(_02118_),
    .A3(_00260_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06795_ (.A1(_00255_),
    .A2(_00259_),
    .B(_00323_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06796_ (.A1(_00263_),
    .A2(_00302_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06797_ (.A1(_00261_),
    .A2(_00303_),
    .B(_00325_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06798_ (.A1(_00289_),
    .A2(_00300_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06799_ (.A1(_00289_),
    .A2(_00300_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06800_ (.A1(_00286_),
    .A2(_00327_),
    .B(_00328_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06801_ (.A1(_02269_),
    .A2(_02802_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06802_ (.A1(_00188_),
    .A2(_00330_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06803_ (.A1(_00290_),
    .A2(_00292_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06804_ (.A1(_00331_),
    .A2(_00332_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06805_ (.A1(_00329_),
    .A2(_00333_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06806_ (.A1(_01749_),
    .A2(_03856_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06807_ (.A1(_00334_),
    .A2(_00335_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06808_ (.A1(_00264_),
    .A2(_00283_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06809_ (.I(_00301_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06810_ (.A1(_00264_),
    .A2(_00283_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06811_ (.A1(_00337_),
    .A2(_00338_),
    .B(_00339_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06812_ (.A1(_00296_),
    .A2(_00299_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06813_ (.A1(_00296_),
    .A2(_00299_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06814_ (.A1(_00293_),
    .A2(_00341_),
    .B(_00342_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06815_ (.A1(_00277_),
    .A2(_00280_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06816_ (.A1(_00275_),
    .A2(_00281_),
    .B(_00344_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06817_ (.A1(net26),
    .A2(_01998_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06818_ (.A1(net25),
    .A2(_02943_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06819_ (.A1(_00330_),
    .A2(_00347_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06820_ (.A1(_00346_),
    .A2(_00348_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06821_ (.A1(_03553_),
    .A2(_03389_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06822_ (.A1(_00295_),
    .A2(_00298_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06823_ (.A1(_00194_),
    .A2(_00350_),
    .B1(_00351_),
    .B2(_00297_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06824_ (.A1(_03629_),
    .A2(_03237_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06825_ (.A1(_02357_),
    .A2(_05628_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06826_ (.A1(_00350_),
    .A2(_00353_),
    .A3(_00354_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06827_ (.A1(_00352_),
    .A2(_00355_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06828_ (.A1(_00349_),
    .A2(_00356_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06829_ (.A1(_00343_),
    .A2(_00345_),
    .A3(_00357_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06830_ (.A1(_00271_),
    .A2(_00282_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06831_ (.A1(_00265_),
    .A2(_00270_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06832_ (.A1(_05359_),
    .A2(_03867_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06833_ (.A1(_02151_),
    .A2(_05413_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06834_ (.A1(net92),
    .A2(net13),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06835_ (.A1(_00265_),
    .A2(_00363_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06836_ (.A1(_00361_),
    .A2(_00362_),
    .B(_00364_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06837_ (.A1(_03640_),
    .A2(_05365_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06838_ (.A1(_02216_),
    .A2(_02889_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06839_ (.A1(net88),
    .A2(_05213_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06840_ (.A1(_00367_),
    .A2(_00368_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06841_ (.A1(_00366_),
    .A2(_00369_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06842_ (.A1(_00360_),
    .A2(_00365_),
    .A3(_00370_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06843_ (.A1(_00273_),
    .A2(_00279_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06844_ (.A1(net86),
    .A2(_02639_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06845_ (.A1(_00177_),
    .A2(_00373_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06846_ (.A1(_00278_),
    .A2(_00372_),
    .B(_00374_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06847_ (.A1(_00268_),
    .A2(_02899_),
    .B1(_01531_),
    .B2(_02226_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06848_ (.A1(_00102_),
    .A2(_00367_),
    .B1(_00376_),
    .B2(_00267_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06849_ (.A1(_02478_),
    .A2(_03356_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06850_ (.A1(_05513_),
    .A2(_00373_),
    .A3(_00378_),
    .Z(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06851_ (.A1(_00377_),
    .A2(_00379_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06852_ (.A1(_00375_),
    .A2(_00380_),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06853_ (.A1(_00371_),
    .A2(_00381_),
    .Z(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06854_ (.A1(_00359_),
    .A2(_00382_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06855_ (.A1(_00358_),
    .A2(_00383_),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06856_ (.A1(_00340_),
    .A2(_00384_),
    .Z(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06857_ (.A1(_00336_),
    .A2(_00385_),
    .Z(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06858_ (.A1(_00326_),
    .A2(_00386_),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06859_ (.A1(_00324_),
    .A2(_00387_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06860_ (.A1(_00322_),
    .A2(_00388_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06861_ (.A1(_00320_),
    .A2(_00389_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06862_ (.A1(_03922_),
    .A2(_00229_),
    .A3(_00239_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06863_ (.A1(_00229_),
    .A2(_00239_),
    .B(_03922_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06864_ (.A1(_05431_),
    .A2(_00392_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06865_ (.I(_05331_),
    .Z(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06866_ (.I(_01401_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06867_ (.I(_03889_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06868_ (.I(_04366_),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06869_ (.A1(_00395_),
    .A2(_00396_),
    .B(_03911_),
    .C(_00397_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06870_ (.A1(_02063_),
    .A2(_00130_),
    .B1(_00394_),
    .B2(_00210_),
    .C(_00398_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06871_ (.A1(_03878_),
    .A2(_05280_),
    .B1(_00396_),
    .B2(_05282_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06872_ (.A1(_00231_),
    .A2(_05180_),
    .B(_00399_),
    .C(_00400_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06873_ (.A1(_00391_),
    .A2(_00393_),
    .B(_00401_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06874_ (.A1(_05446_),
    .A2(_00316_),
    .B1(_00390_),
    .B2(_05496_),
    .C(_00402_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06875_ (.I(_02096_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06876_ (.A1(_00403_),
    .A2(_00396_),
    .A3(_00392_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06877_ (.A1(_00396_),
    .A2(_00392_),
    .B(_00403_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06878_ (.A1(_04097_),
    .A2(_00405_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06879_ (.A1(_00231_),
    .A2(_03933_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06880_ (.A1(_00407_),
    .A2(_00313_),
    .B(_03944_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06881_ (.A1(_00403_),
    .A2(_00408_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06882_ (.A1(_03966_),
    .A2(_02085_),
    .A3(_03955_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06883_ (.A1(_00403_),
    .A2(_03955_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06884_ (.A1(_05444_),
    .A2(_00411_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06885_ (.A1(_05528_),
    .A2(_00409_),
    .B(_00410_),
    .C(_00412_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06886_ (.I(_05384_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06887_ (.A1(_03966_),
    .A2(_00414_),
    .B1(_04269_),
    .B2(_00231_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06888_ (.I(_02063_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06889_ (.I(_02085_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06890_ (.I(_01944_),
    .Z(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06891_ (.A1(_00418_),
    .A2(_00416_),
    .A3(_00417_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06892_ (.A1(_00416_),
    .A2(_00417_),
    .B(_00238_),
    .C(_00419_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06893_ (.I(_00240_),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06894_ (.A1(_03966_),
    .A2(_05380_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06895_ (.A1(_00421_),
    .A2(_00422_),
    .B(_00417_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06896_ (.A1(_00413_),
    .A2(_00415_),
    .A3(_00420_),
    .A4(_00423_),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06897_ (.I(_00244_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06898_ (.A1(_00322_),
    .A2(_00388_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06899_ (.A1(_00322_),
    .A2(_00388_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06900_ (.A1(_00320_),
    .A2(_00426_),
    .B(_00427_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06901_ (.A1(_00326_),
    .A2(_00386_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06902_ (.A1(_00324_),
    .A2(_00387_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06903_ (.A1(_01760_),
    .A2(_03856_),
    .A3(_00334_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06904_ (.A1(_00329_),
    .A2(_00333_),
    .B(_00431_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06905_ (.A1(_00340_),
    .A2(_00384_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06906_ (.A1(_00336_),
    .A2(_00385_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06907_ (.A1(_00433_),
    .A2(_00434_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06908_ (.A1(_00345_),
    .A2(_00357_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06909_ (.A1(_00345_),
    .A2(_00357_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06910_ (.A1(_00343_),
    .A2(_00436_),
    .B(_00437_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06911_ (.A1(_00330_),
    .A2(_00347_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06912_ (.A1(_00346_),
    .A2(_00348_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06913_ (.A1(_00439_),
    .A2(_00440_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06914_ (.A1(_00438_),
    .A2(_00441_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06915_ (.A1(_01760_),
    .A2(_02053_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06916_ (.A1(_00442_),
    .A2(_00443_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06917_ (.A1(_00359_),
    .A2(_00382_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06918_ (.A1(_00358_),
    .A2(_00383_),
    .B(_00445_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06919_ (.A1(_00352_),
    .A2(_00355_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06920_ (.A1(_00349_),
    .A2(_00356_),
    .B(_00447_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06921_ (.A1(_05515_),
    .A2(_00373_),
    .A3(_00378_),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06922_ (.A1(_00377_),
    .A2(_00449_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06923_ (.A1(_00375_),
    .A2(_00380_),
    .B(_00450_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06924_ (.A1(net28),
    .A2(_02020_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06925_ (.A1(net26),
    .A2(_02824_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06926_ (.A1(_00347_),
    .A2(_00453_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06927_ (.A1(_02172_),
    .A2(_02824_),
    .B1(_02965_),
    .B2(net26),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06928_ (.A1(_00454_),
    .A2(_00455_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06929_ (.A1(_00452_),
    .A2(_00456_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06930_ (.A1(_00350_),
    .A2(_00354_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06931_ (.A1(_02357_),
    .A2(_03455_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06932_ (.A1(_00298_),
    .A2(_00459_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06933_ (.A1(_00353_),
    .A2(_00458_),
    .B(_00460_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06934_ (.A1(_02269_),
    .A2(_05324_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06935_ (.A1(_03683_),
    .A2(_05628_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06936_ (.A1(_00459_),
    .A2(_00463_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06937_ (.A1(_00462_),
    .A2(_00464_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06938_ (.A1(_00461_),
    .A2(_00465_),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06939_ (.A1(_00461_),
    .A2(_00465_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06940_ (.A1(_00466_),
    .A2(_00467_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06941_ (.A1(_00457_),
    .A2(_00468_),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06942_ (.A1(_00448_),
    .A2(_00451_),
    .A3(_00469_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06943_ (.A1(_00365_),
    .A2(_00370_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06944_ (.A1(_00365_),
    .A2(_00370_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06945_ (.A1(_00360_),
    .A2(_00471_),
    .A3(_00472_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06946_ (.A1(_00371_),
    .A2(_00381_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06947_ (.A1(_00473_),
    .A2(_00474_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06948_ (.A1(net90),
    .A2(net14),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06949_ (.A1(net12),
    .A2(net93),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06950_ (.A1(_00363_),
    .A2(_00476_),
    .A3(_00477_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06951_ (.A1(_00364_),
    .A2(_00478_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06952_ (.A1(_02216_),
    .A2(_02748_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06953_ (.A1(net87),
    .A2(_02639_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06954_ (.A1(_00268_),
    .A2(_05327_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06955_ (.A1(_00480_),
    .A2(_00481_),
    .A3(_00482_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06956_ (.A1(_00479_),
    .A2(_00483_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06957_ (.A1(_00471_),
    .A2(_00484_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06958_ (.A1(_02401_),
    .A2(net19),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06959_ (.A1(_00373_),
    .A2(_00378_),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06960_ (.A1(_00279_),
    .A2(_00486_),
    .B1(_00487_),
    .B2(_05514_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06961_ (.A1(_00269_),
    .A2(_00480_),
    .B1(_00369_),
    .B2(_00366_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06962_ (.A1(_03553_),
    .A2(_02575_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06963_ (.A1(net85),
    .A2(net20),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06964_ (.A1(_00486_),
    .A2(_00491_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06965_ (.A1(_00490_),
    .A2(_00492_),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06966_ (.A1(_00489_),
    .A2(_00493_),
    .Z(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06967_ (.A1(_00488_),
    .A2(_00494_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06968_ (.A1(_00485_),
    .A2(_00495_),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06969_ (.A1(_00475_),
    .A2(_00496_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06970_ (.A1(_00470_),
    .A2(_00497_),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06971_ (.A1(_00446_),
    .A2(_00498_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06972_ (.A1(_00444_),
    .A2(_00499_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06973_ (.A1(_00432_),
    .A2(_00435_),
    .A3(_00500_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06974_ (.A1(_00429_),
    .A2(_00430_),
    .B(_00501_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06975_ (.A1(_00429_),
    .A2(_00430_),
    .A3(_00501_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06976_ (.A1(_00502_),
    .A2(_00503_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06977_ (.A1(_00428_),
    .A2(_00504_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06978_ (.A1(_00425_),
    .A2(_00505_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06979_ (.A1(_00404_),
    .A2(_00406_),
    .B(_00424_),
    .C(_00506_),
    .ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06980_ (.A1(_00438_),
    .A2(_00441_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06981_ (.A1(_00442_),
    .A2(_00443_),
    .B(_00507_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06982_ (.A1(_00446_),
    .A2(_00498_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06983_ (.I(_00499_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06984_ (.A1(_00444_),
    .A2(_00510_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06985_ (.A1(_00509_),
    .A2(_00511_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06986_ (.A1(_00451_),
    .A2(_00469_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06987_ (.A1(_00451_),
    .A2(_00469_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06988_ (.A1(_00448_),
    .A2(_00513_),
    .B(_00514_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06989_ (.A1(_00452_),
    .A2(_00456_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06990_ (.A1(_00454_),
    .A2(_00516_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06991_ (.A1(_00515_),
    .A2(_00517_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06992_ (.A1(_00475_),
    .A2(_00496_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06993_ (.A1(_00470_),
    .A2(_00497_),
    .B(_00519_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06994_ (.A1(_00471_),
    .A2(_00484_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06995_ (.A1(_00485_),
    .A2(_00495_),
    .B(_00521_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06996_ (.A1(_00364_),
    .A2(_00478_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06997_ (.A1(_00479_),
    .A2(_00483_),
    .B(_00523_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06998_ (.A1(_02074_),
    .A2(_01520_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06999_ (.A1(_00363_),
    .A2(_00477_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07000_ (.A1(_00361_),
    .A2(_00525_),
    .B1(_00526_),
    .B2(_00476_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07001_ (.A1(_02140_),
    .A2(_02748_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07002_ (.A1(_03867_),
    .A2(_05352_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07003_ (.A1(_00525_),
    .A2(_00528_),
    .A3(_00529_),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07004_ (.A1(_00527_),
    .A2(_00530_),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07005_ (.A1(_03651_),
    .A2(_05560_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07006_ (.A1(_02216_),
    .A2(_05327_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07007_ (.A1(_00268_),
    .A2(_05407_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07008_ (.A1(_00533_),
    .A2(_00534_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07009_ (.A1(_00532_),
    .A2(_00535_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07010_ (.A1(_00531_),
    .A2(_00536_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07011_ (.A1(_00524_),
    .A2(_00537_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07012_ (.A1(_02401_),
    .A2(_02532_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07013_ (.A1(_00378_),
    .A2(_00539_),
    .B1(_00492_),
    .B2(_00490_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07014_ (.I(_00540_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07015_ (.A1(_00480_),
    .A2(_00482_),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07016_ (.A1(_00368_),
    .A2(_00533_),
    .B1(_00542_),
    .B2(_00481_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07017_ (.A1(_05524_),
    .A2(_00539_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07018_ (.A1(_02368_),
    .A2(_02586_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07019_ (.A1(_00544_),
    .A2(_00545_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07020_ (.A1(_00543_),
    .A2(_00546_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07021_ (.A1(_00541_),
    .A2(_00547_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07022_ (.A1(_00538_),
    .A2(_00548_),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07023_ (.A1(_00522_),
    .A2(_00549_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07024_ (.I(_00550_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07025_ (.A1(_00457_),
    .A2(_00468_),
    .B(_00466_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07026_ (.A1(_00489_),
    .A2(_00493_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07027_ (.A1(_00488_),
    .A2(_00494_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07028_ (.A1(_00553_),
    .A2(_00554_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07029_ (.A1(net29),
    .A2(_03030_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07030_ (.A1(net28),
    .A2(_02965_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07031_ (.A1(_00453_),
    .A2(_00557_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07032_ (.A1(_00556_),
    .A2(_00558_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07033_ (.A1(_03694_),
    .A2(_03400_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07034_ (.A1(_00354_),
    .A2(_00560_),
    .B1(_00464_),
    .B2(_00462_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07035_ (.A1(_02172_),
    .A2(_05324_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07036_ (.A1(_02269_),
    .A2(_02704_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07037_ (.A1(_00560_),
    .A2(_00563_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07038_ (.A1(_00562_),
    .A2(_00564_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07039_ (.A1(_00561_),
    .A2(_00565_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07040_ (.A1(_00559_),
    .A2(_00566_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07041_ (.A1(_00552_),
    .A2(_00555_),
    .A3(_00567_),
    .Z(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07042_ (.A1(_00551_),
    .A2(_00568_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07043_ (.A1(_00520_),
    .A2(_00569_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07044_ (.A1(_00518_),
    .A2(_00570_),
    .Z(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07045_ (.A1(_00508_),
    .A2(_00512_),
    .A3(_00571_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07046_ (.I(_00435_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07047_ (.A1(_00573_),
    .A2(_00500_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07048_ (.A1(_00573_),
    .A2(_00500_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07049_ (.A1(_00432_),
    .A2(_00574_),
    .B(_00575_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07050_ (.A1(_00572_),
    .A2(_00576_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07051_ (.A1(_00429_),
    .A2(_00430_),
    .A3(_00501_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07052_ (.A1(_00427_),
    .A2(_00502_),
    .B(_00578_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07053_ (.A1(_00319_),
    .A2(_00579_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07054_ (.A1(_00389_),
    .A2(_00502_),
    .A3(_00503_),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07055_ (.A1(_00317_),
    .A2(_00580_),
    .B1(_00581_),
    .B2(_00579_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07056_ (.A1(_00577_),
    .A2(_00582_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07057_ (.I(_05387_),
    .Z(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07058_ (.I(_00584_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07059_ (.A1(_00416_),
    .A2(_00417_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07060_ (.A1(_00586_),
    .A2(_00405_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07061_ (.I(_00234_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07062_ (.A1(_00416_),
    .A2(_00585_),
    .B1(_00587_),
    .B2(_05317_),
    .C(_00588_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07063_ (.A1(_05115_),
    .A2(_00583_),
    .B(_00589_),
    .ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07064_ (.A1(_00572_),
    .A2(_00576_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07065_ (.A1(_00317_),
    .A2(_00580_),
    .B1(_00581_),
    .B2(_00579_),
    .C(_00577_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07066_ (.A1(_00590_),
    .A2(_00591_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07067_ (.A1(_00515_),
    .A2(_00517_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07068_ (.A1(_00520_),
    .A2(_00569_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07069_ (.A1(_00518_),
    .A2(_00570_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07070_ (.A1(_00594_),
    .A2(_00595_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07071_ (.I(_00555_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07072_ (.A1(_00597_),
    .A2(_00567_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07073_ (.A1(_00597_),
    .A2(_00567_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07074_ (.A1(_00552_),
    .A2(_00598_),
    .B(_00599_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07075_ (.A1(_00453_),
    .A2(_00557_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07076_ (.A1(_00556_),
    .A2(_00558_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07077_ (.A1(_00601_),
    .A2(_00602_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07078_ (.A1(_00600_),
    .A2(_00603_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07079_ (.A1(_00522_),
    .A2(_00549_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07080_ (.A1(_00551_),
    .A2(_00568_),
    .B(_00605_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07081_ (.A1(_00524_),
    .A2(_00537_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07082_ (.A1(_00538_),
    .A2(_00548_),
    .B(_00607_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07083_ (.I(_00527_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07084_ (.A1(_00531_),
    .A2(_00536_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07085_ (.A1(_00609_),
    .A2(_00530_),
    .B(_00610_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07086_ (.A1(_02074_),
    .A2(_02889_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07087_ (.A1(_00525_),
    .A2(_00529_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07088_ (.A1(_00363_),
    .A2(_00612_),
    .B1(_00613_),
    .B2(_00528_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07089_ (.A1(_02140_),
    .A2(_05365_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07090_ (.A1(net92),
    .A2(_02748_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07091_ (.A1(_00612_),
    .A2(_00616_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07092_ (.A1(_00615_),
    .A2(_00617_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07093_ (.A1(_00614_),
    .A2(_00618_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07094_ (.A1(_03651_),
    .A2(_02543_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07095_ (.A1(_02226_),
    .A2(_03367_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07096_ (.A1(_00534_),
    .A2(_00621_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07097_ (.A1(_02324_),
    .A2(_05560_),
    .B1(_05408_),
    .B2(_02237_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07098_ (.A1(_00622_),
    .A2(_00623_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07099_ (.A1(_00620_),
    .A2(_00624_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07100_ (.A1(_00619_),
    .A2(_00625_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07101_ (.I(_00626_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07102_ (.A1(_00611_),
    .A2(_00627_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07103_ (.I(_00628_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07104_ (.A1(_02423_),
    .A2(_03564_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07105_ (.A1(_00491_),
    .A2(_00630_),
    .B1(_00544_),
    .B2(_00545_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07106_ (.A1(_00533_),
    .A2(_00534_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07107_ (.A1(_00532_),
    .A2(_00535_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07108_ (.A1(_00632_),
    .A2(_00633_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07109_ (.A1(_03694_),
    .A2(_02596_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07110_ (.A1(_02368_),
    .A2(_02489_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07111_ (.A1(_00630_),
    .A2(_00636_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07112_ (.A1(_00635_),
    .A2(_00637_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07113_ (.A1(_00634_),
    .A2(_00638_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07114_ (.A1(_00631_),
    .A2(_00639_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07115_ (.A1(_00629_),
    .A2(_00640_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07116_ (.A1(_00608_),
    .A2(_00641_),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07117_ (.A1(_00561_),
    .A2(_00565_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07118_ (.A1(_00559_),
    .A2(_00566_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07119_ (.A1(_00643_),
    .A2(_00644_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07120_ (.I(_00645_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07121_ (.A1(_00543_),
    .A2(_00546_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07122_ (.A1(_00541_),
    .A2(_00547_),
    .B(_00647_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07123_ (.A1(net28),
    .A2(_02845_),
    .B1(_04539_),
    .B2(_02053_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07124_ (.A1(_02053_),
    .A2(_02845_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07125_ (.A1(_00557_),
    .A2(_00650_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07126_ (.A1(_00649_),
    .A2(_00651_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07127_ (.A1(_02280_),
    .A2(_03411_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07128_ (.A1(_00463_),
    .A2(_00653_),
    .B1(_00564_),
    .B2(_00562_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07129_ (.A1(_02107_),
    .A2(_05325_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07130_ (.A1(_02183_),
    .A2(_02715_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07131_ (.A1(_00653_),
    .A2(_00656_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07132_ (.A1(_00655_),
    .A2(_00657_),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07133_ (.A1(_00654_),
    .A2(_00658_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07134_ (.A1(_00652_),
    .A2(_00659_),
    .Z(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07135_ (.A1(_00646_),
    .A2(_00648_),
    .A3(_00660_),
    .Z(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07136_ (.A1(_00642_),
    .A2(_00661_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07137_ (.A1(_00606_),
    .A2(_00662_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07138_ (.A1(_00604_),
    .A2(_00663_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07139_ (.A1(_00593_),
    .A2(_00596_),
    .A3(_00664_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07140_ (.A1(_00512_),
    .A2(_00571_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07141_ (.A1(_00512_),
    .A2(_00571_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07142_ (.A1(_00508_),
    .A2(_00666_),
    .B(_00667_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07143_ (.A1(_00665_),
    .A2(_00668_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07144_ (.A1(_00592_),
    .A2(_00669_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07145_ (.I(_05665_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07146_ (.A1(_00592_),
    .A2(_00669_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07147_ (.A1(_00671_),
    .A2(_00672_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07148_ (.I(_01249_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07149_ (.A1(_00670_),
    .A2(_00673_),
    .B(_00674_),
    .ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07150_ (.I(_05344_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07151_ (.I(_00668_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07152_ (.A1(_00665_),
    .A2(_00676_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07153_ (.A1(_00592_),
    .A2(_00669_),
    .B(_00677_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07154_ (.A1(_00594_),
    .A2(_00595_),
    .A3(_00664_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07155_ (.A1(_00594_),
    .A2(_00595_),
    .B(_00664_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07156_ (.A1(_00593_),
    .A2(_00679_),
    .B(_00680_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07157_ (.A1(_00606_),
    .A2(_00662_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07158_ (.A1(_00604_),
    .A2(_00663_),
    .B(_00682_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07159_ (.I(_00639_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07160_ (.A1(_00631_),
    .A2(_00684_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07161_ (.A1(_00634_),
    .A2(_00638_),
    .B(_00685_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07162_ (.A1(_02183_),
    .A2(_03509_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07163_ (.A1(_00563_),
    .A2(_00687_),
    .B1(_00657_),
    .B2(_00655_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07164_ (.A1(_03900_),
    .A2(_05325_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07165_ (.A1(_00650_),
    .A2(_00687_),
    .A3(_00689_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07166_ (.A1(_00686_),
    .A2(_00688_),
    .A3(_00690_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07167_ (.A1(_00600_),
    .A2(_00603_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07168_ (.A1(_03705_),
    .A2(_02607_),
    .A3(_00637_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07169_ (.A1(_05584_),
    .A2(_00693_),
    .B(_05651_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07170_ (.A1(_05652_),
    .A2(_00693_),
    .B(_00694_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07171_ (.A1(_00692_),
    .A2(_00695_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07172_ (.I(_00608_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07173_ (.A1(_00697_),
    .A2(_00641_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07174_ (.A1(_00642_),
    .A2(_00661_),
    .B(_00698_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07175_ (.A1(_00648_),
    .A2(_00660_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07176_ (.A1(_00648_),
    .A2(_00660_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07177_ (.A1(_00646_),
    .A2(_00700_),
    .B(_00701_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07178_ (.A1(_03694_),
    .A2(_02500_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07179_ (.A1(_02151_),
    .A2(_02661_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07180_ (.A1(_03867_),
    .A2(_03204_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07181_ (.A1(_02324_),
    .A2(_02553_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07182_ (.A1(_00704_),
    .A2(_00705_),
    .A3(_00706_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07183_ (.A1(_00621_),
    .A2(_00703_),
    .A3(_00707_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07184_ (.A1(_00534_),
    .A2(_00621_),
    .B1(_00624_),
    .B2(_00620_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07185_ (.A1(_02074_),
    .A2(_02780_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07186_ (.A1(_00529_),
    .A2(_00710_),
    .B1(_00617_),
    .B2(_00615_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07187_ (.A1(_00708_),
    .A2(_00709_),
    .A3(_00711_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07188_ (.A1(_00611_),
    .A2(_00627_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07189_ (.A1(_00629_),
    .A2(_00640_),
    .B(_00713_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07190_ (.A1(_00614_),
    .A2(_00618_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07191_ (.A1(_00619_),
    .A2(_00625_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07192_ (.A1(_00715_),
    .A2(_00716_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07193_ (.A1(_03716_),
    .A2(_03574_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07194_ (.A1(_02280_),
    .A2(_02596_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07195_ (.A1(_00710_),
    .A2(_00718_),
    .A3(_00719_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07196_ (.A1(_00714_),
    .A2(_00717_),
    .A3(_00720_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07197_ (.A1(_00654_),
    .A2(_00658_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07198_ (.A1(_00652_),
    .A2(_00659_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07199_ (.A1(_00722_),
    .A2(_00723_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07200_ (.A1(_02107_),
    .A2(_02726_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07201_ (.A1(_00724_),
    .A2(_00725_),
    .Z(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07202_ (.A1(_00712_),
    .A2(_00721_),
    .A3(_00726_),
    .Z(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07203_ (.A1(_00651_),
    .A2(_00702_),
    .A3(_00727_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07204_ (.A1(_00696_),
    .A2(_00699_),
    .A3(_00728_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07205_ (.A1(_00691_),
    .A2(_00729_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07206_ (.A1(_00681_),
    .A2(_00683_),
    .A3(_00730_),
    .Z(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07207_ (.A1(_00678_),
    .A2(_00731_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07208_ (.A1(_00678_),
    .A2(_00731_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07209_ (.I(_04626_),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07210_ (.I(_00734_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07211_ (.A1(_00675_),
    .A2(_00732_),
    .A3(_00733_),
    .B(_00735_),
    .ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07212_ (.I(net5),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07213_ (.I(_00736_),
    .Z(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07214_ (.I(_00737_),
    .Z(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07215_ (.I(_00738_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07216_ (.I(_00739_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07217_ (.I(_00740_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07218_ (.I(_00739_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07219_ (.I(net69),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07220_ (.I(_00743_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07221_ (.A1(_00742_),
    .A2(_00744_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07222_ (.I(net69),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07223_ (.A1(_00740_),
    .A2(_00746_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07224_ (.A1(_00745_),
    .A2(_00747_),
    .B(_01498_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07225_ (.I(net16),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07226_ (.I(_00749_),
    .Z(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07227_ (.I(_00750_),
    .Z(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07228_ (.I(_00751_),
    .Z(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07229_ (.I(_00752_),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07230_ (.I(_00753_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07231_ (.I(_00744_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07232_ (.I(_00755_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07233_ (.I(_00756_),
    .Z(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07234_ (.I(_00757_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07235_ (.A1(_00758_),
    .A2(_01890_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07236_ (.A1(_01825_),
    .A2(_00759_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _07237_ (.A1(_00754_),
    .A2(_01662_),
    .B1(_01738_),
    .B2(_00758_),
    .C1(_00741_),
    .C2(_00760_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07238_ (.A1(_00741_),
    .A2(_01249_),
    .B(_00748_),
    .C(_00761_),
    .ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07239_ (.I(_04919_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07240_ (.I(_00752_),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07241_ (.I(net80),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07242_ (.I(_00764_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07243_ (.I(_00765_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07244_ (.I(_00766_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07245_ (.I(_00767_),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07246_ (.A1(_00763_),
    .A2(_00768_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07247_ (.I(net11),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07248_ (.I(_00770_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07249_ (.I(net75),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07250_ (.A1(_00771_),
    .A2(_00772_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07251_ (.I(net9),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07252_ (.I(_00774_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07253_ (.I(_00775_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07254_ (.I(net73),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07255_ (.I(_00777_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07256_ (.A1(_00776_),
    .A2(_00778_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07257_ (.I(net8),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07258_ (.I(_00780_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07259_ (.I(_00781_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07260_ (.I(_00782_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07261_ (.I(net72),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07262_ (.I(_00784_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07263_ (.I(_00785_),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07264_ (.I(_00786_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07265_ (.A1(_00783_),
    .A2(_00787_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07266_ (.I(net7),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07267_ (.I(_00789_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07268_ (.I(_00790_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07269_ (.I(net71),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07270_ (.I(_00792_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07271_ (.I(_00793_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07272_ (.A1(_00791_),
    .A2(_00794_),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07273_ (.I(net68),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07274_ (.I(net132),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07275_ (.I(_00797_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07276_ (.I(_00798_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07277_ (.I(_00799_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07278_ (.A1(_00796_),
    .A2(_00800_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07279_ (.A1(_00796_),
    .A2(_00799_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07280_ (.I(net67),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07281_ (.I(_00803_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07282_ (.I(net131),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07283_ (.I(_00805_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07284_ (.I(_00806_),
    .Z(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07285_ (.A1(_00804_),
    .A2(_00807_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07286_ (.I(net66),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07287_ (.I(_00809_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07288_ (.I(_00810_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07289_ (.I(_00811_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07290_ (.I(net130),
    .Z(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07291_ (.I(_00813_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07292_ (.I(_00814_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07293_ (.I(_00815_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07294_ (.I(_00816_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07295_ (.A1(_00812_),
    .A2(_00817_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07296_ (.I(net60),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07297_ (.I(_00819_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07298_ (.I(_00820_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07299_ (.I(_00821_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07300_ (.I(net124),
    .Z(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07301_ (.I(_00823_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07302_ (.I(_00824_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07303_ (.I(_00825_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07304_ (.A1(_00822_),
    .A2(_00826_),
    .Z(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07305_ (.I(net38),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07306_ (.I(_00828_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07307_ (.I(_00829_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07308_ (.I(_00830_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07309_ (.I(_00831_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07310_ (.I(net102),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07311_ (.I(_00833_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07312_ (.I(_00834_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07313_ (.I(_00835_),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07314_ (.I(_00836_),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07315_ (.I(_00837_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07316_ (.A1(_00832_),
    .A2(_00838_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07317_ (.I(_00839_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07318_ (.A1(_00831_),
    .A2(_00836_),
    .Z(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07319_ (.A1(_00830_),
    .A2(_00835_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07320_ (.I(_00842_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07321_ (.I(net27),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07322_ (.I(_00844_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07323_ (.I(_00845_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07324_ (.I(_00846_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07325_ (.I(net91),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07326_ (.I(_00848_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07327_ (.I(_00849_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07328_ (.I(_00850_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07329_ (.I(_00851_),
    .Z(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07330_ (.I(_00852_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07331_ (.A1(_00847_),
    .A2(_00853_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07332_ (.I(_00763_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07333_ (.A1(_00855_),
    .A2(_00768_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07334_ (.A1(_00742_),
    .A2(_00744_),
    .B(_00769_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07335_ (.A1(_00846_),
    .A2(_00849_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07336_ (.I(_00858_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07337_ (.A1(_00847_),
    .A2(_00852_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07338_ (.A1(_00859_),
    .A2(_00860_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07339_ (.A1(_00856_),
    .A2(_00857_),
    .B(_00861_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07340_ (.A1(_00841_),
    .A2(_00843_),
    .B1(_00854_),
    .B2(_00862_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07341_ (.A1(_00841_),
    .A2(_00843_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07342_ (.I(_00768_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07343_ (.A1(_00855_),
    .A2(_00865_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07344_ (.A1(_00745_),
    .A2(_00769_),
    .B(_00866_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07345_ (.A1(_00864_),
    .A2(_00861_),
    .A3(_00867_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07346_ (.A1(_00840_),
    .A2(_00863_),
    .B(_00868_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07347_ (.I(net49),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07348_ (.I(_00870_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07349_ (.I(_00871_),
    .Z(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07350_ (.I(_00872_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07351_ (.I(net113),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07352_ (.I(_00874_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07353_ (.A1(_00873_),
    .A2(_00875_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07354_ (.I(net113),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07355_ (.A1(_00871_),
    .A2(_00877_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07356_ (.A1(_00876_),
    .A2(_00878_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07357_ (.A1(_00821_),
    .A2(_00826_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07358_ (.I(_00872_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07359_ (.A1(_00881_),
    .A2(_00875_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07360_ (.A1(_00869_),
    .A2(_00879_),
    .B(_00880_),
    .C(_00882_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07361_ (.I(net65),
    .Z(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07362_ (.I(_00884_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07363_ (.I(_00885_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07364_ (.I(_00886_),
    .Z(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07365_ (.I(net129),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07366_ (.I(_00888_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07367_ (.I(_00889_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07368_ (.A1(_00887_),
    .A2(_00890_),
    .Z(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07369_ (.I(net65),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07370_ (.I(_00892_),
    .Z(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07371_ (.I(net129),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07372_ (.I(_00894_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07373_ (.A1(_00893_),
    .A2(_00895_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07374_ (.A1(_00891_),
    .A2(_00896_),
    .Z(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07375_ (.I(_00887_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07376_ (.I(_00890_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07377_ (.A1(_00898_),
    .A2(_00899_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07378_ (.A1(_00827_),
    .A2(_00883_),
    .A3(_00897_),
    .B(_00900_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07379_ (.A1(_00812_),
    .A2(_00817_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07380_ (.I(net67),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07381_ (.I(_00903_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07382_ (.I(_00904_),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07383_ (.I(net131),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07384_ (.I(_00906_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07385_ (.A1(_00905_),
    .A2(_00907_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07386_ (.A1(_00818_),
    .A2(_00901_),
    .B(_00902_),
    .C(_00908_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07387_ (.A1(_00802_),
    .A2(_00808_),
    .A3(_00909_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07388_ (.I(net6),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07389_ (.I(_00911_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07390_ (.I(net70),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07391_ (.I(_00913_),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07392_ (.I(_00914_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07393_ (.I(_00915_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07394_ (.A1(_00912_),
    .A2(_00916_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07395_ (.I(net6),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07396_ (.I(_00918_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07397_ (.I(_00919_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07398_ (.I(_00914_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07399_ (.A1(_00920_),
    .A2(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07400_ (.A1(_00917_),
    .A2(_00922_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07401_ (.A1(_00912_),
    .A2(_00921_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07402_ (.A1(_00801_),
    .A2(_00910_),
    .A3(_00923_),
    .B(_00924_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07403_ (.A1(_00791_),
    .A2(_00794_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07404_ (.A1(_00783_),
    .A2(_00786_),
    .B1(_00795_),
    .B2(_00925_),
    .C(_00926_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07405_ (.I(_00778_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07406_ (.A1(_00776_),
    .A2(_00928_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07407_ (.A1(_00779_),
    .A2(_00788_),
    .A3(_00927_),
    .B(_00929_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07408_ (.I(net10),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07409_ (.I(_00931_),
    .Z(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07410_ (.I(net74),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07411_ (.I(_00933_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07412_ (.I(_00934_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07413_ (.A1(_00932_),
    .A2(_00935_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07414_ (.A1(_00932_),
    .A2(_00935_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07415_ (.A1(_00930_),
    .A2(_00936_),
    .B(_00937_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07416_ (.I(_00771_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07417_ (.I(_00772_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07418_ (.A1(_00939_),
    .A2(_00940_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07419_ (.A1(_00773_),
    .A2(_00938_),
    .B(_00941_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07420_ (.I(_00942_),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07421_ (.I(_00943_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07422_ (.I(_00944_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07423_ (.I(_00943_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07424_ (.A1(_00742_),
    .A2(_00758_),
    .B(_00946_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07425_ (.A1(_00747_),
    .A2(_00945_),
    .B(_00947_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07426_ (.A1(_00769_),
    .A2(_00948_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07427_ (.I(_05497_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07428_ (.I(_01836_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07429_ (.A1(_00758_),
    .A2(_00754_),
    .B1(_00865_),
    .B2(_00741_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07430_ (.I(_00743_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07431_ (.I(_00953_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07432_ (.A1(_00740_),
    .A2(_00954_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07433_ (.A1(_00753_),
    .A2(_00768_),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07434_ (.I(_00956_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07435_ (.A1(_00955_),
    .A2(_00957_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07436_ (.I(_05591_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07437_ (.A1(_00951_),
    .A2(_00952_),
    .A3(_00958_),
    .B1(_00959_),
    .B2(_00957_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07438_ (.A1(_00865_),
    .A2(_00950_),
    .B(_00960_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07439_ (.A1(_00740_),
    .A2(_00756_),
    .A3(_00769_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07440_ (.A1(_00855_),
    .A2(_00865_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07441_ (.I(_01412_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07442_ (.A1(_00955_),
    .A2(_00963_),
    .B(_00964_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07443_ (.I(_04626_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07444_ (.I(_00847_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07445_ (.I(_05506_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07446_ (.A1(_00967_),
    .A2(_04637_),
    .B1(_00968_),
    .B2(_00741_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07447_ (.A1(_00754_),
    .A2(_00966_),
    .B1(_00963_),
    .B2(_04388_),
    .C(_00969_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07448_ (.A1(_00962_),
    .A2(_00965_),
    .B(_00970_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07449_ (.A1(_00762_),
    .A2(_00949_),
    .B(_00961_),
    .C(_00971_),
    .ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07450_ (.I(_00861_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07451_ (.A1(_00856_),
    .A2(_00857_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07452_ (.I(_00944_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07453_ (.A1(_00867_),
    .A2(_00946_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07454_ (.A1(_00973_),
    .A2(_00974_),
    .B(_00975_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07455_ (.A1(_00972_),
    .A2(_00976_),
    .B(_05291_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07456_ (.A1(_00972_),
    .A2(_00976_),
    .B(_00977_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07457_ (.I(_01423_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07458_ (.A1(_00957_),
    .A2(_00972_),
    .A3(_00962_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07459_ (.A1(_00957_),
    .A2(_00962_),
    .B(_00861_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07460_ (.A1(_00979_),
    .A2(_00980_),
    .A3(_00981_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07461_ (.I(_01640_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07462_ (.I(_05387_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07463_ (.I(_00859_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07464_ (.A1(_05202_),
    .A2(_00985_),
    .B(_00860_),
    .C(_04377_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07465_ (.A1(_00832_),
    .A2(_00983_),
    .B1(_00984_),
    .B2(_00754_),
    .C(_00986_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07466_ (.I(_04150_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07467_ (.I(_04204_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07468_ (.A1(_00852_),
    .A2(_00988_),
    .B1(_00985_),
    .B2(_00989_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07469_ (.A1(_00967_),
    .A2(_00734_),
    .B(_00987_),
    .C(_00990_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07470_ (.I(_01847_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07471_ (.A1(_00739_),
    .A2(_00851_),
    .A3(_00763_),
    .A4(_00767_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07472_ (.A1(_00738_),
    .A2(_00851_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07473_ (.A1(_00956_),
    .A2(_00994_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07474_ (.A1(_00993_),
    .A2(_00995_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07475_ (.A1(_00953_),
    .A2(_00847_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07476_ (.A1(_00996_),
    .A2(_00997_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07477_ (.I(_00998_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07478_ (.A1(_00996_),
    .A2(_00997_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07479_ (.A1(_00958_),
    .A2(_00999_),
    .A3(_01000_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07480_ (.A1(_00999_),
    .A2(_01000_),
    .B(_00958_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07481_ (.A1(_00992_),
    .A2(_01001_),
    .A3(_01002_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _07482_ (.A1(_00978_),
    .A2(_00982_),
    .A3(_00991_),
    .A4(_01003_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07483_ (.I(_01004_),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07484_ (.A1(_00967_),
    .A2(_00853_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07485_ (.A1(_00972_),
    .A2(_00867_),
    .B(_01005_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07486_ (.I(_00943_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07487_ (.I(_01007_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07488_ (.A1(_00854_),
    .A2(_00862_),
    .A3(_01008_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07489_ (.A1(_00945_),
    .A2(_01006_),
    .B(_01009_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07490_ (.A1(_00864_),
    .A2(_01010_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07491_ (.A1(_00864_),
    .A2(_01010_),
    .B(_05663_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07492_ (.A1(_00851_),
    .A2(_00763_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07493_ (.A1(_00846_),
    .A2(_00767_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07494_ (.A1(_00739_),
    .A2(_00836_),
    .ZN(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07495_ (.A1(_01013_),
    .A2(_01014_),
    .A3(_01015_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07496_ (.A1(_00743_),
    .A2(_00831_),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07497_ (.A1(_00993_),
    .A2(_01017_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07498_ (.A1(_01016_),
    .A2(_01018_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07499_ (.A1(_00998_),
    .A2(_01019_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07500_ (.I(_00999_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07501_ (.I(_01019_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07502_ (.A1(_01021_),
    .A2(_01001_),
    .A3(_01022_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07503_ (.A1(_01001_),
    .A2(_01022_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07504_ (.A1(_01020_),
    .A2(_01023_),
    .A3(_01024_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07505_ (.A1(_00985_),
    .A2(_00981_),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07506_ (.A1(_00864_),
    .A2(_01026_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07507_ (.I(_04086_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07508_ (.I(net38),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07509_ (.I(_01029_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07510_ (.A1(_01030_),
    .A2(_00833_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07511_ (.A1(_01944_),
    .A2(_01031_),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07512_ (.A1(_01346_),
    .A2(_00841_),
    .A3(_01032_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07513_ (.A1(_00881_),
    .A2(_00211_),
    .B1(_00212_),
    .B2(_00967_),
    .C(_01033_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07514_ (.I(_04193_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07515_ (.A1(_00837_),
    .A2(_00217_),
    .B1(_01031_),
    .B2(_01035_),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07516_ (.A1(_00832_),
    .A2(_04290_),
    .B(_01034_),
    .C(_01036_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07517_ (.A1(_05666_),
    .A2(_01025_),
    .B1(_01027_),
    .B2(_01028_),
    .C(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07518_ (.A1(_01011_),
    .A2(_01012_),
    .B(_01038_),
    .ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07519_ (.I(_00879_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07520_ (.I(_01039_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07521_ (.A1(_00840_),
    .A2(_00863_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07522_ (.I0(_01041_),
    .I1(_00869_),
    .S(_00974_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07523_ (.A1(_01040_),
    .A2(_01042_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07524_ (.A1(_01040_),
    .A2(_01042_),
    .B(_05663_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07525_ (.A1(_00993_),
    .A2(_01017_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07526_ (.A1(_01016_),
    .A2(_01018_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07527_ (.A1(_01045_),
    .A2(_01046_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07528_ (.I(_00736_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07529_ (.I(_01048_),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07530_ (.I(_00877_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07531_ (.A1(_01049_),
    .A2(_01050_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07532_ (.A1(_00834_),
    .A2(_00751_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07533_ (.A1(_00830_),
    .A2(_00766_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07534_ (.A1(_00858_),
    .A2(_01052_),
    .A3(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07535_ (.A1(_01051_),
    .A2(_01054_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07536_ (.A1(_00738_),
    .A2(_00835_),
    .B1(_00850_),
    .B2(_00752_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07537_ (.A1(_00994_),
    .A2(_01052_),
    .B1(_01056_),
    .B2(_01014_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07538_ (.A1(net69),
    .A2(_00871_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07539_ (.A1(_01057_),
    .A2(_01058_),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07540_ (.A1(_01055_),
    .A2(_01059_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07541_ (.A1(_01047_),
    .A2(_01060_),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07542_ (.A1(_01020_),
    .A2(_01061_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07543_ (.A1(_01024_),
    .A2(_01062_),
    .Z(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07544_ (.A1(_00985_),
    .A2(_00981_),
    .B(_00841_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07545_ (.A1(_00843_),
    .A2(_01040_),
    .A3(_01064_),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07546_ (.A1(_00843_),
    .A2(_01064_),
    .B(_01039_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07547_ (.A1(_01065_),
    .A2(_01066_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07548_ (.I(_00822_),
    .Z(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07549_ (.A1(_00881_),
    .A2(_00049_),
    .B1(_01368_),
    .B2(_01040_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07550_ (.A1(_01068_),
    .A2(_05435_),
    .B1(_00876_),
    .B2(_05437_),
    .C(_01069_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07551_ (.I(_01050_),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07552_ (.I(_01071_),
    .Z(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07553_ (.I(_05506_),
    .Z(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07554_ (.I(net49),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07555_ (.A1(_01074_),
    .A2(_00874_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07556_ (.A1(_01072_),
    .A2(_05326_),
    .B1(_01073_),
    .B2(_00832_),
    .C1(_01075_),
    .C2(_05512_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07557_ (.A1(_01070_),
    .A2(_01076_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07558_ (.A1(_05666_),
    .A2(_01063_),
    .B1(_01067_),
    .B2(_01028_),
    .C(_01077_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07559_ (.A1(_01043_),
    .A2(_01044_),
    .B(_01078_),
    .ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07560_ (.A1(_00999_),
    .A2(_01019_),
    .A3(_01061_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07561_ (.A1(_01024_),
    .A2(_01062_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07562_ (.A1(_01045_),
    .A2(_01046_),
    .B(_01060_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07563_ (.A1(_00755_),
    .A2(_00872_),
    .A3(_01057_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07564_ (.A1(_01055_),
    .A2(_01059_),
    .B(_01082_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07565_ (.A1(_00836_),
    .A2(_00753_),
    .B(_00859_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07566_ (.I(net102),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07567_ (.I(_01085_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07568_ (.I(net27),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07569_ (.I(_01088_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07570_ (.A1(_01087_),
    .A2(_01089_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07571_ (.A1(_01053_),
    .A2(_01084_),
    .B1(_01090_),
    .B2(_01013_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07572_ (.A1(_00743_),
    .A2(_00821_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07573_ (.A1(_01091_),
    .A2(_01092_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07574_ (.A1(_01051_),
    .A2(_01054_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07575_ (.I(net124),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07576_ (.I(_01095_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07577_ (.A1(_01048_),
    .A2(_01096_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07578_ (.A1(_01071_),
    .A2(_00752_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07579_ (.A1(_01049_),
    .A2(_00824_),
    .A3(_01050_),
    .A4(_00751_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07580_ (.A1(_01098_),
    .A2(_01099_),
    .B(_01100_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07581_ (.I(_01074_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07582_ (.A1(_01102_),
    .A2(_00764_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07583_ (.A1(_00830_),
    .A2(_00849_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07584_ (.A1(_01090_),
    .A2(_01103_),
    .A3(_01104_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07585_ (.A1(_01101_),
    .A2(_01105_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07586_ (.A1(_01094_),
    .A2(_01106_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07587_ (.A1(_01093_),
    .A2(_01107_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07588_ (.A1(_01083_),
    .A2(_01109_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07589_ (.A1(_01081_),
    .A2(_01110_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07590_ (.A1(_01079_),
    .A2(_01080_),
    .A3(_01111_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07591_ (.I(_05665_),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07592_ (.A1(_01079_),
    .A2(_01080_),
    .B(_01111_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07593_ (.A1(_01113_),
    .A2(_01114_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07594_ (.A1(_00827_),
    .A2(_00880_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07595_ (.A1(_01075_),
    .A2(_01066_),
    .B(_01116_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07596_ (.I(_01423_),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07597_ (.I(_01116_),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07598_ (.A1(_01075_),
    .A2(_01066_),
    .A3(_01120_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07599_ (.A1(_01118_),
    .A2(_01121_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07600_ (.I(_01803_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07601_ (.A1(_00887_),
    .A2(_04323_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07602_ (.A1(_01068_),
    .A2(_05169_),
    .B(_01124_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07603_ (.A1(_00881_),
    .A2(_00584_),
    .B1(_01120_),
    .B2(_01123_),
    .C(_01125_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07604_ (.A1(_00819_),
    .A2(_01095_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07605_ (.I(_01127_),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07606_ (.A1(_01879_),
    .A2(_01128_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07607_ (.A1(_01068_),
    .A2(_05320_),
    .B1(_00988_),
    .B2(_00825_),
    .C(_01129_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07608_ (.A1(_01126_),
    .A2(_01131_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07609_ (.A1(_01117_),
    .A2(_01122_),
    .B(_01132_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07610_ (.A1(_00873_),
    .A2(_01072_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07611_ (.A1(_01041_),
    .A2(_01039_),
    .B(_01134_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07612_ (.A1(_00869_),
    .A2(_01039_),
    .B(_00882_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07613_ (.I(_00942_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07614_ (.I0(_01135_),
    .I1(_01136_),
    .S(_01137_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07615_ (.I(_05444_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07616_ (.A1(_01120_),
    .A2(_01138_),
    .B(_01139_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07617_ (.A1(_01120_),
    .A2(_01138_),
    .B(_01140_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07618_ (.A1(_01112_),
    .A2(_01115_),
    .B(_01133_),
    .C(_01142_),
    .ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07619_ (.A1(_00891_),
    .A2(_00896_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07620_ (.I(_01143_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07621_ (.A1(_00822_),
    .A2(_00826_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07622_ (.A1(_00880_),
    .A2(_01135_),
    .B(_01145_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07623_ (.A1(_01008_),
    .A2(_01146_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07624_ (.A1(_00827_),
    .A2(_00883_),
    .A3(_01008_),
    .B(_01147_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07625_ (.A1(_01144_),
    .A2(_01148_),
    .Z(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07626_ (.A1(_01144_),
    .A2(_01148_),
    .B(_05663_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07627_ (.I(_05294_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07628_ (.A1(_01081_),
    .A2(_01110_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07629_ (.A1(_01083_),
    .A2(_01109_),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07630_ (.A1(_01101_),
    .A2(_01105_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07631_ (.I(net60),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07632_ (.I(_01156_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07633_ (.A1(_01157_),
    .A2(_00764_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07634_ (.A1(_00871_),
    .A2(_00848_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07635_ (.A1(_01031_),
    .A2(_01158_),
    .A3(_01159_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07636_ (.I(_00749_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07637_ (.A1(_01096_),
    .A2(_01161_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07638_ (.A1(_00877_),
    .A2(_00845_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07639_ (.A1(_00737_),
    .A2(_00889_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07640_ (.A1(_01163_),
    .A2(_01164_),
    .A3(_01165_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07641_ (.A1(_01100_),
    .A2(_01160_),
    .A3(_01166_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07642_ (.A1(_01155_),
    .A2(_01167_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07643_ (.I(_01168_),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07644_ (.A1(_01094_),
    .A2(_01106_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07645_ (.A1(net69),
    .A2(_00886_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07646_ (.A1(_01090_),
    .A2(_01104_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07647_ (.A1(_01031_),
    .A2(_00859_),
    .B1(_01103_),
    .B2(_01172_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07648_ (.A1(_01170_),
    .A2(_01171_),
    .A3(_01174_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07649_ (.A1(_01169_),
    .A2(_01175_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07650_ (.A1(_00755_),
    .A2(_00821_),
    .A3(_01091_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07651_ (.A1(_01093_),
    .A2(_01107_),
    .B(_01177_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07652_ (.A1(_01176_),
    .A2(_01178_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07653_ (.A1(_01154_),
    .A2(_01179_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07654_ (.A1(_01153_),
    .A2(_01114_),
    .A3(_01180_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07655_ (.A1(_01153_),
    .A2(_01114_),
    .B(_01180_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07656_ (.A1(_01181_),
    .A2(_01182_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07657_ (.A1(_01144_),
    .A2(_01117_),
    .A3(_01128_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07658_ (.A1(_01117_),
    .A2(_01128_),
    .B(_01144_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07659_ (.A1(_00045_),
    .A2(_01186_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07660_ (.I(_00812_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07661_ (.I(_05519_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07662_ (.A1(_01188_),
    .A2(_04334_),
    .B1(_01189_),
    .B2(_00897_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07663_ (.A1(_00884_),
    .A2(_00894_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07664_ (.I(_04193_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07665_ (.I(_01192_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07666_ (.A1(_00899_),
    .A2(_04161_),
    .B1(_01191_),
    .B2(_01193_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07667_ (.A1(_00898_),
    .A2(_00131_),
    .B1(_00394_),
    .B2(_01068_),
    .C1(_00891_),
    .C2(_05586_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07668_ (.A1(_01190_),
    .A2(_01194_),
    .A3(_01196_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07669_ (.A1(_01152_),
    .A2(_01183_),
    .B1(_01185_),
    .B2(_01187_),
    .C(_01197_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07670_ (.A1(_01149_),
    .A2(_01150_),
    .B(_01198_),
    .ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07671_ (.I(_01188_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07672_ (.A1(_01199_),
    .A2(_00816_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07673_ (.A1(_01200_),
    .A2(_00902_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07674_ (.A1(_00898_),
    .A2(_00899_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07675_ (.A1(_01143_),
    .A2(_01146_),
    .B(_01202_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07676_ (.A1(_01007_),
    .A2(_01203_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07677_ (.A1(_00901_),
    .A2(_01007_),
    .B(_01204_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07678_ (.A1(_01201_),
    .A2(_01206_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07679_ (.A1(_01154_),
    .A2(_01179_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07680_ (.A1(_01176_),
    .A2(_01178_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07681_ (.A1(_01169_),
    .A2(_01175_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07682_ (.A1(_01170_),
    .A2(_01174_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07683_ (.A1(_01170_),
    .A2(_01174_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07684_ (.A1(_01171_),
    .A2(_01211_),
    .B(_01212_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07685_ (.A1(_01049_),
    .A2(_00814_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07686_ (.A1(_01051_),
    .A2(_01163_),
    .Z(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07687_ (.A1(_01215_),
    .A2(_01166_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07688_ (.A1(_01215_),
    .A2(_01166_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07689_ (.A1(_01160_),
    .A2(_01217_),
    .B(_01218_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07690_ (.I(_01219_),
    .Z(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07691_ (.A1(_00885_),
    .A2(_00765_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07692_ (.A1(_00870_),
    .A2(_00833_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07693_ (.I(net91),
    .Z(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07694_ (.A1(_00819_),
    .A2(_01223_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07695_ (.A1(_01222_),
    .A2(_01224_),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07696_ (.A1(_01221_),
    .A2(_01225_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07697_ (.A1(net129),
    .A2(net16),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07698_ (.A1(_00736_),
    .A2(_00888_),
    .B1(_00823_),
    .B2(_01161_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07699_ (.A1(_01098_),
    .A2(_01228_),
    .B1(_01229_),
    .B2(_01164_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07700_ (.A1(net113),
    .A2(_01029_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07701_ (.A1(_01095_),
    .A2(_00844_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07702_ (.A1(_01228_),
    .A2(_01231_),
    .A3(_01232_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07703_ (.A1(_01230_),
    .A2(_01233_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07704_ (.A1(_01226_),
    .A2(_01234_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07705_ (.I(_01235_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07706_ (.A1(_01214_),
    .A2(_01220_),
    .A3(_01236_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07707_ (.A1(_00953_),
    .A2(_00812_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07708_ (.A1(_01155_),
    .A2(_01167_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07709_ (.A1(_00842_),
    .A2(_01159_),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07710_ (.A1(_01158_),
    .A2(_01241_),
    .B1(_01222_),
    .B2(_01104_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07711_ (.A1(_01240_),
    .A2(_01242_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07712_ (.A1(_01237_),
    .A2(_01239_),
    .A3(_01243_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07713_ (.A1(_01210_),
    .A2(_01213_),
    .A3(_01244_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07714_ (.A1(_01209_),
    .A2(_01245_),
    .Z(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07715_ (.A1(_01208_),
    .A2(_01182_),
    .A3(_01246_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07716_ (.A1(_01208_),
    .A2(_01182_),
    .B(_01246_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07717_ (.A1(_05295_),
    .A2(_01247_),
    .A3(_01248_),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07718_ (.I(_05497_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07719_ (.A1(_01191_),
    .A2(_01186_),
    .A3(_01201_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07720_ (.A1(_01191_),
    .A2(_01186_),
    .B(_01201_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07721_ (.A1(_01252_),
    .A2(_01253_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07722_ (.I(_05502_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07723_ (.I(_00905_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07724_ (.I(_05504_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07725_ (.A1(_01256_),
    .A2(_00983_),
    .B1(_01257_),
    .B2(_01199_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07726_ (.A1(net66),
    .A2(net130),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07727_ (.I(_01259_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07728_ (.I(_01261_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07729_ (.I(_01192_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07730_ (.A1(_00887_),
    .A2(_00984_),
    .B1(_01262_),
    .B2(_01263_),
    .ZN(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07731_ (.I(_05436_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07732_ (.A1(_01188_),
    .A2(_01265_),
    .B1(_01189_),
    .B2(_01201_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07733_ (.A1(_01258_),
    .A2(_01264_),
    .A3(_01266_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07734_ (.A1(_00816_),
    .A2(_01251_),
    .B1(_01254_),
    .B2(_01255_),
    .C(_01267_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07735_ (.A1(_00762_),
    .A2(_01207_),
    .B(_01250_),
    .C(_01268_),
    .ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07736_ (.A1(_00804_),
    .A2(_00907_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07737_ (.A1(_01256_),
    .A2(_00807_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07738_ (.A1(_01269_),
    .A2(_01271_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07739_ (.I(_01272_),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07740_ (.A1(_00902_),
    .A2(_01203_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07741_ (.A1(_00818_),
    .A2(_00901_),
    .B(_01137_),
    .C(_00902_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07742_ (.A1(_00818_),
    .A2(_00945_),
    .A3(_01274_),
    .B(_01275_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07743_ (.A1(_01273_),
    .A2(_01276_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07744_ (.A1(_01273_),
    .A2(_01276_),
    .B(_01976_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07745_ (.A1(_01209_),
    .A2(_01245_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07746_ (.I(_01279_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07747_ (.A1(_01210_),
    .A2(_01244_),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07748_ (.A1(_01210_),
    .A2(_01244_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07749_ (.A1(_01213_),
    .A2(_01282_),
    .B(_01283_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07750_ (.A1(_01239_),
    .A2(_01243_),
    .Z(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07751_ (.A1(_01237_),
    .A2(_01285_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07752_ (.A1(_01239_),
    .A2(_01243_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07753_ (.A1(_01240_),
    .A2(_01242_),
    .B(_01287_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07754_ (.A1(_01219_),
    .A2(_01235_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07755_ (.A1(_01220_),
    .A2(_01236_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07756_ (.A1(_01214_),
    .A2(_01289_),
    .A3(_01290_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07757_ (.A1(_00746_),
    .A2(_00804_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07758_ (.A1(_01222_),
    .A2(_01224_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07759_ (.A1(_01221_),
    .A2(_01225_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07760_ (.A1(_01294_),
    .A2(_01295_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07761_ (.A1(_01289_),
    .A2(_01293_),
    .A3(_01296_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07762_ (.A1(_01049_),
    .A2(_00806_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07763_ (.A1(_00815_),
    .A2(_00753_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07764_ (.A1(_00805_),
    .A2(_00749_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07765_ (.A1(_01214_),
    .A2(_01300_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07766_ (.A1(_01298_),
    .A2(_01299_),
    .B(_01301_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07767_ (.A1(_01230_),
    .A2(_01233_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07768_ (.A1(_01226_),
    .A2(_01234_),
    .B(_01304_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07769_ (.A1(_00811_),
    .A2(_00765_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07770_ (.A1(_00893_),
    .A2(_01157_),
    .A3(_01087_),
    .A4(_00848_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07771_ (.A1(_00820_),
    .A2(_00834_),
    .B1(_00848_),
    .B2(_00885_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07772_ (.A1(_01307_),
    .A2(_01308_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07773_ (.A1(_01306_),
    .A2(_01309_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07774_ (.A1(_00894_),
    .A2(_01088_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07775_ (.A1(_00824_),
    .A2(_00846_),
    .B1(_00751_),
    .B2(_00889_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07776_ (.A1(_01163_),
    .A2(_01311_),
    .B1(_01312_),
    .B2(_01231_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07777_ (.A1(_00823_),
    .A2(_01030_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07778_ (.A1(_01075_),
    .A2(_01311_),
    .A3(_01315_),
    .Z(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07779_ (.A1(_01313_),
    .A2(_01316_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07780_ (.A1(_01310_),
    .A2(_01317_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07781_ (.A1(_01305_),
    .A2(_01318_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07782_ (.A1(_01302_),
    .A2(_01319_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07783_ (.A1(_01291_),
    .A2(_01297_),
    .A3(_01320_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07784_ (.A1(_01286_),
    .A2(_01288_),
    .A3(_01321_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07785_ (.A1(_01284_),
    .A2(_01322_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07786_ (.I(_01323_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07787_ (.A1(_01280_),
    .A2(_01248_),
    .A3(_01324_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07788_ (.A1(_01280_),
    .A2(_01248_),
    .B(_01324_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07789_ (.A1(_05344_),
    .A2(_01327_),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07790_ (.A1(_01326_),
    .A2(_01328_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07791_ (.A1(_01253_),
    .A2(_01261_),
    .A3(_01273_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07792_ (.A1(_01253_),
    .A2(_01261_),
    .B(_01272_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07793_ (.A1(_00979_),
    .A2(_01331_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07794_ (.I(net68),
    .Z(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07795_ (.I(_01333_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07796_ (.I(_01334_),
    .Z(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07797_ (.I(_01335_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07798_ (.I(_04323_),
    .Z(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07799_ (.A1(_01256_),
    .A2(_05169_),
    .B1(_01379_),
    .B2(_01273_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07800_ (.A1(_01337_),
    .A2(_01338_),
    .B1(_01269_),
    .B2(_00237_),
    .C(_01339_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07801_ (.A1(_00803_),
    .A2(_00907_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07802_ (.A1(_00807_),
    .A2(_04161_),
    .B1(_00584_),
    .B2(_01188_),
    .C1(_01341_),
    .C2(_01193_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07803_ (.A1(_01340_),
    .A2(_01342_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07804_ (.A1(_01330_),
    .A2(_01332_),
    .B(_01343_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07805_ (.A1(_01277_),
    .A2(_01278_),
    .B(_01329_),
    .C(_01344_),
    .ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07806_ (.I(_05445_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07807_ (.A1(_01337_),
    .A2(_00800_),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07808_ (.A1(_01269_),
    .A2(_01271_),
    .Z(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07809_ (.A1(_00818_),
    .A2(_01348_),
    .A3(_01274_),
    .B(_00908_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07810_ (.A1(_00808_),
    .A2(_00909_),
    .A3(_00944_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07811_ (.A1(_01137_),
    .A2(_01349_),
    .B(_01350_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07812_ (.A1(_01347_),
    .A2(_01351_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07813_ (.A1(_01284_),
    .A2(_01322_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07814_ (.A1(_01353_),
    .A2(_01327_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07815_ (.A1(_01237_),
    .A2(_01285_),
    .A3(_01321_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07816_ (.A1(_01286_),
    .A2(_01321_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07817_ (.A1(_01288_),
    .A2(_01356_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07818_ (.A1(_01220_),
    .A2(_01236_),
    .B(_01296_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07819_ (.A1(_01220_),
    .A2(_01236_),
    .A3(_01296_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07820_ (.A1(_01293_),
    .A2(_01359_),
    .B(_01360_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07821_ (.I(_01361_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07822_ (.A1(_01291_),
    .A2(_01320_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07823_ (.A1(_01291_),
    .A2(_01320_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07824_ (.A1(_01297_),
    .A2(_01363_),
    .B(_01364_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07825_ (.A1(_01302_),
    .A2(_01319_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07826_ (.A1(_00813_),
    .A2(_01088_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07827_ (.A1(_00737_),
    .A2(_00799_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07828_ (.A1(_01300_),
    .A2(_01367_),
    .A3(_01369_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07829_ (.A1(_01301_),
    .A2(_01370_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07830_ (.A1(_01313_),
    .A2(_01316_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07831_ (.A1(_01310_),
    .A2(_01317_),
    .B(_01372_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07832_ (.A1(_00884_),
    .A2(_01087_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07833_ (.I(net80),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07834_ (.A1(_00804_),
    .A2(_01375_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07835_ (.A1(_00810_),
    .A2(_00849_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07836_ (.A1(_01374_),
    .A2(_01376_),
    .A3(_01377_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07837_ (.A1(net129),
    .A2(_00828_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07838_ (.I(_01095_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07839_ (.A1(_01381_),
    .A2(_00829_),
    .B1(_00845_),
    .B2(_00895_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07840_ (.A1(_01232_),
    .A2(_01380_),
    .B1(_01382_),
    .B2(_00878_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07841_ (.A1(_01156_),
    .A2(net113),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07842_ (.A1(net124),
    .A2(_01074_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07843_ (.A1(_01380_),
    .A2(_01384_),
    .A3(_01385_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07844_ (.A1(_01383_),
    .A2(_01386_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07845_ (.A1(_01378_),
    .A2(_01387_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07846_ (.A1(_01373_),
    .A2(_01388_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07847_ (.A1(_01371_),
    .A2(_01389_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07848_ (.A1(_01366_),
    .A2(_01391_),
    .Z(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07849_ (.A1(_00953_),
    .A2(_01335_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07850_ (.A1(_01305_),
    .A2(_01318_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07851_ (.A1(_01306_),
    .A2(_01309_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07852_ (.A1(_01307_),
    .A2(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07853_ (.A1(_01394_),
    .A2(_01396_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07854_ (.A1(_01393_),
    .A2(_01397_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07855_ (.A1(_01392_),
    .A2(_01398_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07856_ (.A1(_01362_),
    .A2(_01365_),
    .A3(_01399_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07857_ (.A1(_01355_),
    .A2(_01358_),
    .B(_01400_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07858_ (.A1(_01355_),
    .A2(_01358_),
    .A3(_01400_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07859_ (.A1(_01402_),
    .A2(_01403_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07860_ (.A1(_01354_),
    .A2(_01404_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07861_ (.I(_05104_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07862_ (.A1(_01341_),
    .A2(_01331_),
    .A3(_01347_),
    .Z(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07863_ (.A1(_01341_),
    .A2(_01331_),
    .B(_01347_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07864_ (.A1(_01407_),
    .A2(_01408_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07865_ (.I(_05506_),
    .Z(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07866_ (.A1(_01335_),
    .A2(_00800_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07867_ (.I(_01411_),
    .Z(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07868_ (.A1(_01879_),
    .A2(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07869_ (.A1(_01256_),
    .A2(_01410_),
    .B(_01414_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07870_ (.I(_00920_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07871_ (.I(_05510_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07872_ (.I(_05504_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07873_ (.A1(_01416_),
    .A2(_01417_),
    .B1(_01418_),
    .B2(_00796_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07874_ (.A1(_01337_),
    .A2(_05517_),
    .B1(_00133_),
    .B2(_01347_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07875_ (.A1(_01415_),
    .A2(_01419_),
    .A3(_01420_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07876_ (.A1(_00800_),
    .A2(_05644_),
    .B1(_01409_),
    .B2(_05648_),
    .C(_01421_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07877_ (.A1(_01345_),
    .A2(_01352_),
    .B1(_01405_),
    .B2(_01406_),
    .C(_01422_),
    .ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07878_ (.A1(_00801_),
    .A2(_00910_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07879_ (.A1(_00802_),
    .A2(_01349_),
    .B(_00801_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07880_ (.A1(_00974_),
    .A2(_01425_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07881_ (.A1(_01424_),
    .A2(_00945_),
    .B(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07882_ (.A1(_00923_),
    .A2(_01427_),
    .B(_05445_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07883_ (.A1(_00923_),
    .A2(_01427_),
    .B(_01428_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07884_ (.I(_05665_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07885_ (.A1(_01365_),
    .A2(_01399_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07886_ (.A1(_01365_),
    .A2(_01399_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07887_ (.A1(_01362_),
    .A2(_01431_),
    .B(_01432_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07888_ (.A1(_01307_),
    .A2(_01395_),
    .B(_01394_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07889_ (.A1(_01393_),
    .A2(_01397_),
    .B(_01435_),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07890_ (.A1(_01302_),
    .A2(_01319_),
    .A3(_01391_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07891_ (.A1(_01392_),
    .A2(_01398_),
    .B(_01437_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07892_ (.A1(_01371_),
    .A2(_01389_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07893_ (.A1(_00736_),
    .A2(_00913_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07894_ (.A1(_00798_),
    .A2(_00750_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07895_ (.A1(_01300_),
    .A2(_01369_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07896_ (.A1(_01298_),
    .A2(_01441_),
    .B1(_01442_),
    .B2(_01367_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07897_ (.A1(_00813_),
    .A2(_00829_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07898_ (.A1(_00806_),
    .A2(_01089_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07899_ (.A1(_01441_),
    .A2(_01445_),
    .A3(_01446_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07900_ (.A1(_01443_),
    .A2(_01447_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07901_ (.A1(_01440_),
    .A2(_01448_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07902_ (.A1(_01383_),
    .A2(_01386_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07903_ (.A1(_01378_),
    .A2(_01387_),
    .B(_01450_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07904_ (.A1(_01301_),
    .A2(_01370_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07905_ (.A1(net66),
    .A2(_01085_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07906_ (.A1(_00796_),
    .A2(_01375_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07907_ (.A1(_00903_),
    .A2(net91),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07908_ (.A1(_01453_),
    .A2(_01454_),
    .A3(_01456_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07909_ (.A1(_00894_),
    .A2(net49),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07910_ (.A1(_01380_),
    .A2(_01385_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _07911_ (.A1(_01315_),
    .A2(_01458_),
    .B1(_01459_),
    .B2(_01384_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07912_ (.A1(_00884_),
    .A2(_00877_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07913_ (.A1(_01127_),
    .A2(_01458_),
    .A3(_01461_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07914_ (.A1(_01457_),
    .A2(_01460_),
    .A3(_01462_),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07915_ (.A1(_01452_),
    .A2(_01463_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07916_ (.A1(_01451_),
    .A2(_01464_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07917_ (.A1(_01449_),
    .A2(_01465_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07918_ (.A1(_00744_),
    .A2(_00919_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07919_ (.A1(_01373_),
    .A2(_01388_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07920_ (.A1(_01374_),
    .A2(_01377_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07921_ (.A1(_01374_),
    .A2(_01377_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07922_ (.A1(_01376_),
    .A2(_01470_),
    .B(_01471_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07923_ (.A1(_01469_),
    .A2(_01472_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07924_ (.A1(_01468_),
    .A2(_01473_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07925_ (.A1(_01439_),
    .A2(_01467_),
    .A3(_01474_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07926_ (.A1(_01438_),
    .A2(_01475_),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07927_ (.A1(_01436_),
    .A2(_01476_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07928_ (.A1(_01434_),
    .A2(_01478_),
    .Z(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07929_ (.I(_01479_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07930_ (.I(_01402_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07931_ (.A1(_01353_),
    .A2(_01327_),
    .A3(_01481_),
    .B(_01403_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07932_ (.A1(_01480_),
    .A2(_01482_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07933_ (.A1(_00917_),
    .A2(_00922_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07934_ (.A1(_01484_),
    .A2(_01408_),
    .A3(_01413_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07935_ (.A1(_01408_),
    .A2(_01413_),
    .B(_01484_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07936_ (.A1(_00979_),
    .A2(_01486_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07937_ (.I(_00791_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07938_ (.I(_01489_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07939_ (.A1(_01416_),
    .A2(_05169_),
    .B1(_01379_),
    .B2(_01484_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07940_ (.A1(_01490_),
    .A2(_01338_),
    .B1(_00917_),
    .B2(_00237_),
    .C(_01491_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07941_ (.I(_04150_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07942_ (.A1(_00912_),
    .A2(_00916_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07943_ (.A1(_00921_),
    .A2(_01493_),
    .B1(_00984_),
    .B2(_01337_),
    .C1(_01494_),
    .C2(_01263_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07944_ (.A1(_01492_),
    .A2(_01495_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07945_ (.A1(_01430_),
    .A2(_01483_),
    .B1(_01485_),
    .B2(_01487_),
    .C(_01496_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07946_ (.A1(_01429_),
    .A2(_01497_),
    .ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07947_ (.I(_01489_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07948_ (.I(_00793_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07949_ (.A1(_01499_),
    .A2(_01500_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07950_ (.A1(_00795_),
    .A2(_01501_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07951_ (.A1(_01416_),
    .A2(_00916_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07952_ (.A1(_00920_),
    .A2(_00916_),
    .B1(_00802_),
    .B2(_01349_),
    .C(_00801_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07953_ (.A1(_01503_),
    .A2(_00943_),
    .A3(_01504_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07954_ (.A1(_00925_),
    .A2(_00946_),
    .B(_01505_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07955_ (.A1(_01502_),
    .A2(_01506_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07956_ (.A1(_01434_),
    .A2(_01478_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07957_ (.A1(_01480_),
    .A2(_01482_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07958_ (.A1(_01508_),
    .A2(_01510_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07959_ (.A1(_01438_),
    .A2(_01475_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07960_ (.A1(_01436_),
    .A2(_01476_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07961_ (.A1(_01512_),
    .A2(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07962_ (.A1(_01469_),
    .A2(_01472_),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07963_ (.A1(_01468_),
    .A2(_01473_),
    .B(_01515_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07964_ (.A1(_01439_),
    .A2(_01467_),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07965_ (.A1(_01439_),
    .A2(_01467_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07966_ (.A1(_01517_),
    .A2(_01474_),
    .B(_01518_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07967_ (.A1(_00954_),
    .A2(_00791_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07968_ (.A1(_01452_),
    .A2(_01463_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07969_ (.A1(_01451_),
    .A2(_01464_),
    .B(_01522_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07970_ (.A1(_01453_),
    .A2(_01456_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07971_ (.A1(_00903_),
    .A2(_01085_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07972_ (.A1(_01377_),
    .A2(_01525_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07973_ (.A1(_01454_),
    .A2(_01524_),
    .B(_01526_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07974_ (.A1(_01523_),
    .A2(_01527_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07975_ (.A1(_01521_),
    .A2(_01528_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07976_ (.A1(_01449_),
    .A2(_01465_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07977_ (.A1(_01440_),
    .A2(_01448_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07978_ (.A1(_01460_),
    .A2(_01462_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07979_ (.A1(_01460_),
    .A2(_01462_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07980_ (.A1(_01457_),
    .A2(_01533_),
    .B(_01534_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07981_ (.A1(_01443_),
    .A2(_01447_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07982_ (.A1(_00911_),
    .A2(_01375_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07983_ (.A1(_01333_),
    .A2(_01223_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07984_ (.A1(_01525_),
    .A2(_01537_),
    .A3(_01538_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07985_ (.A1(_01127_),
    .A2(_01458_),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07986_ (.A1(_00888_),
    .A2(_01157_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _07987_ (.A1(_01461_),
    .A2(_01540_),
    .B1(_01541_),
    .B2(_01385_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07988_ (.A1(_00809_),
    .A2(_00874_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07989_ (.A1(_00893_),
    .A2(_01096_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07990_ (.A1(_01541_),
    .A2(_01544_),
    .A3(_01545_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07991_ (.A1(_01539_),
    .A2(_01543_),
    .A3(_01546_),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07992_ (.A1(_01536_),
    .A2(_01547_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07993_ (.A1(_01535_),
    .A2(_01548_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07994_ (.A1(_00737_),
    .A2(_00792_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07995_ (.A1(_00915_),
    .A2(_00855_),
    .B(_01550_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07996_ (.A1(_00792_),
    .A2(_00750_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07997_ (.A1(_01440_),
    .A2(_01552_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07998_ (.I(_01554_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07999_ (.A1(_01551_),
    .A2(_01555_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08000_ (.A1(_00798_),
    .A2(_01089_),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08001_ (.A1(_01441_),
    .A2(_01446_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08002_ (.A1(_01300_),
    .A2(_01557_),
    .B1(_01558_),
    .B2(_01445_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08003_ (.A1(_00814_),
    .A2(_01102_),
    .ZN(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08004_ (.A1(_00805_),
    .A2(_00829_),
    .ZN(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08005_ (.A1(_01557_),
    .A2(_01560_),
    .A3(_01561_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08006_ (.A1(_01559_),
    .A2(_01562_),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08007_ (.A1(_01556_),
    .A2(_01563_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08008_ (.A1(_01532_),
    .A2(_01549_),
    .A3(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08009_ (.A1(_01530_),
    .A2(_01566_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08010_ (.A1(_01529_),
    .A2(_01567_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08011_ (.A1(_01516_),
    .A2(_01519_),
    .A3(_01568_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08012_ (.A1(_01514_),
    .A2(_01569_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08013_ (.A1(_01511_),
    .A2(_01570_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08014_ (.A1(_01494_),
    .A2(_01486_),
    .A3(_01502_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08015_ (.A1(_01494_),
    .A2(_01486_),
    .B(_01502_),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08016_ (.A1(_01572_),
    .A2(_01573_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08017_ (.A1(_01416_),
    .A2(_00126_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08018_ (.I(_05281_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08019_ (.A1(_01490_),
    .A2(_01500_),
    .A3(_01577_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08020_ (.I(_00782_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08021_ (.A1(_01579_),
    .A2(_00211_),
    .B1(_00131_),
    .B2(_01499_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08022_ (.A1(_01490_),
    .A2(_05319_),
    .B1(_05519_),
    .B2(_01502_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08023_ (.A1(_01576_),
    .A2(_01578_),
    .A3(_01580_),
    .A4(_01581_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08024_ (.A1(_01500_),
    .A2(_05644_),
    .B1(_01574_),
    .B2(_05648_),
    .C(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08025_ (.A1(_01345_),
    .A2(_01507_),
    .B1(_01571_),
    .B2(_01406_),
    .C(_01583_),
    .ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08026_ (.A1(_00782_),
    .A2(_00787_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08027_ (.A1(_01579_),
    .A2(_00787_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08028_ (.A1(_01584_),
    .A2(_01586_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08029_ (.I(_01587_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08030_ (.A1(_00926_),
    .A2(_01503_),
    .A3(_01504_),
    .B(_00795_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08031_ (.A1(_00795_),
    .A2(_00925_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08032_ (.A1(_01501_),
    .A2(_01590_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08033_ (.I0(_01589_),
    .I1(_01591_),
    .S(_00974_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08034_ (.A1(_01588_),
    .A2(_01592_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08035_ (.A1(_01588_),
    .A2(_01592_),
    .B(_01976_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08036_ (.A1(_01512_),
    .A2(_01513_),
    .B(_01569_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08037_ (.A1(_01512_),
    .A2(_01513_),
    .A3(_01569_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08038_ (.A1(_01508_),
    .A2(_01595_),
    .B(_01597_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08039_ (.A1(_01480_),
    .A2(_01482_),
    .A3(_01570_),
    .B(_01598_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08040_ (.A1(_01519_),
    .A2(_01568_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08041_ (.A1(_01519_),
    .A2(_01568_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08042_ (.A1(_01516_),
    .A2(_01600_),
    .B(_01601_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08043_ (.A1(_00757_),
    .A2(_01489_),
    .A3(_01528_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08044_ (.A1(_01523_),
    .A2(_01527_),
    .B(_01603_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08045_ (.A1(_01449_),
    .A2(_01465_),
    .A3(_01566_),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08046_ (.A1(_01529_),
    .A2(_01567_),
    .B(_01605_),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08047_ (.A1(_00954_),
    .A2(_00781_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08048_ (.A1(_01536_),
    .A2(_01547_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08049_ (.A1(_01535_),
    .A2(_01548_),
    .B(_01609_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08050_ (.A1(_01525_),
    .A2(_01538_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08051_ (.A1(_01333_),
    .A2(_01085_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08052_ (.A1(_01456_),
    .A2(_01612_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08053_ (.A1(_01537_),
    .A2(_01611_),
    .B(_01613_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08054_ (.A1(_01610_),
    .A2(_01614_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08055_ (.A1(_01608_),
    .A2(_01615_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08056_ (.A1(_01532_),
    .A2(_01565_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08057_ (.A1(_01532_),
    .A2(_01565_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08058_ (.A1(_01549_),
    .A2(_01617_),
    .B(_01619_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08059_ (.A1(_01551_),
    .A2(_01555_),
    .A3(_01563_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08060_ (.A1(_00913_),
    .A2(_01089_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08061_ (.A1(_00738_),
    .A2(_00786_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08062_ (.A1(_01552_),
    .A2(_01622_),
    .A3(_01623_),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08063_ (.A1(net132),
    .A2(_01029_),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08064_ (.A1(_01557_),
    .A2(_01561_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08065_ (.A1(_01446_),
    .A2(_01625_),
    .B1(_01626_),
    .B2(_01560_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08066_ (.A1(net130),
    .A2(net60),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08067_ (.A1(_00906_),
    .A2(_01074_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08068_ (.A1(_01625_),
    .A2(_01628_),
    .A3(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08069_ (.A1(_01554_),
    .A2(_01631_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08070_ (.A1(_01627_),
    .A2(_01632_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08071_ (.A1(_01624_),
    .A2(_01633_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08072_ (.A1(_01621_),
    .A2(_01634_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08073_ (.A1(_01543_),
    .A2(_01546_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08074_ (.A1(_01543_),
    .A2(_01546_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08075_ (.A1(_01539_),
    .A2(_01636_),
    .B(_01637_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08076_ (.A1(_01559_),
    .A2(_01562_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08077_ (.A1(net7),
    .A2(_00764_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08078_ (.A1(net6),
    .A2(net91),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08079_ (.A1(_01612_),
    .A2(_01641_),
    .A3(_01642_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08080_ (.I(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08081_ (.A1(_00895_),
    .A2(_00820_),
    .B1(_01381_),
    .B2(_00893_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08082_ (.A1(_00896_),
    .A2(_01128_),
    .B1(_01544_),
    .B2(_01645_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08083_ (.A1(_00904_),
    .A2(_00874_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08084_ (.A1(_00810_),
    .A2(_01381_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08085_ (.A1(_01191_),
    .A2(_01647_),
    .A3(_01648_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08086_ (.A1(_01644_),
    .A2(_01646_),
    .A3(_01649_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08087_ (.A1(_01639_),
    .A2(_01650_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08088_ (.A1(_01638_),
    .A2(_01652_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08089_ (.A1(_01635_),
    .A2(_01653_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08090_ (.A1(_01620_),
    .A2(_01654_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08091_ (.A1(_01616_),
    .A2(_01655_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08092_ (.A1(_01606_),
    .A2(_01656_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08093_ (.A1(_01604_),
    .A2(_01657_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08094_ (.A1(_01602_),
    .A2(_01658_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08095_ (.A1(_01599_),
    .A2(_01659_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08096_ (.A1(_01489_),
    .A2(_01500_),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08097_ (.A1(_01588_),
    .A2(_01573_),
    .A3(_01661_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08098_ (.A1(_01573_),
    .A2(_01661_),
    .B(_01587_),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08099_ (.A1(_01663_),
    .A2(_01664_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08100_ (.I(_00775_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08101_ (.I(_01584_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08102_ (.A1(_00395_),
    .A2(_01667_),
    .B(_01586_),
    .C(_00397_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08103_ (.A1(_01666_),
    .A2(_05191_),
    .B1(_05267_),
    .B2(_01490_),
    .C(_01668_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08104_ (.A1(_00787_),
    .A2(_00217_),
    .B1(_01667_),
    .B2(_01035_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08105_ (.A1(_01579_),
    .A2(_01238_),
    .B(_01669_),
    .C(_01670_),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08106_ (.A1(_01152_),
    .A2(_01660_),
    .B1(_01665_),
    .B2(_01028_),
    .C(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08107_ (.A1(_01593_),
    .A2(_01594_),
    .B(_01672_),
    .ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08108_ (.A1(_00776_),
    .A2(_00928_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08109_ (.A1(_00779_),
    .A2(_01674_),
    .Z(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08110_ (.A1(_01588_),
    .A2(_01589_),
    .B(_00788_),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08111_ (.A1(_00788_),
    .A2(_00927_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08112_ (.I0(_01676_),
    .I1(_01677_),
    .S(_00944_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08113_ (.A1(_01675_),
    .A2(_01678_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08114_ (.A1(_01667_),
    .A2(_01664_),
    .B(_01675_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08115_ (.A1(_01667_),
    .A2(_01664_),
    .A3(_01675_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08116_ (.A1(_00964_),
    .A2(_01681_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08117_ (.A1(_00776_),
    .A2(_00234_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08118_ (.I(_00932_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08119_ (.A1(_01685_),
    .A2(_01651_),
    .B1(_00126_),
    .B2(_01579_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08120_ (.A1(_01666_),
    .A2(_01265_),
    .B1(_01675_),
    .B2(_01123_),
    .ZN(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08121_ (.A1(_01666_),
    .A2(_00928_),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08122_ (.A1(_01879_),
    .A2(_01688_),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08123_ (.A1(_00928_),
    .A2(_04161_),
    .B(_01689_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08124_ (.A1(_01684_),
    .A2(_01686_),
    .A3(_01687_),
    .A4(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08125_ (.A1(_01602_),
    .A2(_01658_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08126_ (.A1(_01599_),
    .A2(_01659_),
    .B(_01692_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08127_ (.A1(_01606_),
    .A2(_01656_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08128_ (.A1(_01604_),
    .A2(_01657_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08129_ (.A1(_00757_),
    .A2(_00782_),
    .A3(_01615_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08130_ (.A1(_01610_),
    .A2(_01614_),
    .B(_01697_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08131_ (.A1(_01620_),
    .A2(_01654_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08132_ (.A1(_01616_),
    .A2(_01655_),
    .B(_01699_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08133_ (.A1(_00954_),
    .A2(_00774_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08134_ (.A1(_01639_),
    .A2(_01650_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08135_ (.A1(_01638_),
    .A2(_01652_),
    .B(_01702_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08136_ (.A1(_01612_),
    .A2(_01642_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08137_ (.A1(_00918_),
    .A2(_00833_),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08138_ (.A1(_01538_),
    .A2(_01706_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08139_ (.A1(_01641_),
    .A2(_01704_),
    .B(_01707_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08140_ (.A1(_01703_),
    .A2(_01708_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08141_ (.A1(_01701_),
    .A2(_01709_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08142_ (.A1(_01551_),
    .A2(_01555_),
    .A3(_01563_),
    .A4(_01634_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08143_ (.A1(_01635_),
    .A2(_01653_),
    .B(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08144_ (.A1(_01624_),
    .A2(_01633_),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08145_ (.A1(net5),
    .A2(_00777_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08146_ (.A1(net72),
    .A2(net16),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08147_ (.A1(net70),
    .A2(_01029_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08148_ (.I(net71),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08149_ (.A1(_01718_),
    .A2(_00844_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08150_ (.A1(_01715_),
    .A2(_01717_),
    .A3(_01719_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08151_ (.A1(_01714_),
    .A2(_01720_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08152_ (.A1(_01625_),
    .A2(_01630_),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08153_ (.A1(_00797_),
    .A2(net49),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08154_ (.A1(_01561_),
    .A2(_01723_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08155_ (.A1(_01628_),
    .A2(_01722_),
    .B(_01724_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08156_ (.A1(_01048_),
    .A2(_00785_),
    .B1(_00792_),
    .B2(_01161_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08157_ (.A1(_01550_),
    .A2(_01715_),
    .B1(_01726_),
    .B2(_01622_),
    .ZN(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08158_ (.A1(net130),
    .A2(_00892_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08159_ (.A1(_00805_),
    .A2(_01157_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08160_ (.A1(_01723_),
    .A2(_01729_),
    .A3(_01730_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08161_ (.A1(_01728_),
    .A2(_01731_),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08162_ (.A1(_01725_),
    .A2(_01732_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08163_ (.A1(_01721_),
    .A2(_01733_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08164_ (.A1(_01646_),
    .A2(_01649_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08165_ (.A1(_01646_),
    .A2(_01649_),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08166_ (.A1(_01644_),
    .A2(_01735_),
    .B(_01736_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08167_ (.A1(_01555_),
    .A2(_01631_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08168_ (.A1(_01554_),
    .A2(_01631_),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08169_ (.A1(_01627_),
    .A2(_01739_),
    .B(_01740_),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08170_ (.A1(_00780_),
    .A2(_00765_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08171_ (.A1(_00789_),
    .A2(_01223_),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08172_ (.A1(_01706_),
    .A2(_01743_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08173_ (.A1(_01742_),
    .A2(_01744_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08174_ (.A1(_00896_),
    .A2(_01648_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08175_ (.A1(_00810_),
    .A2(_00889_),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08176_ (.A1(_01647_),
    .A2(_01746_),
    .B1(_01747_),
    .B2(_01545_),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08177_ (.A1(_01334_),
    .A2(_01050_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08178_ (.A1(_00904_),
    .A2(_01381_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08179_ (.A1(_01747_),
    .A2(_01750_),
    .A3(_01751_),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08180_ (.A1(_01745_),
    .A2(_01748_),
    .A3(_01752_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08181_ (.A1(_01737_),
    .A2(_01741_),
    .A3(_01753_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08182_ (.A1(_01713_),
    .A2(_01734_),
    .A3(_01754_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08183_ (.A1(_01712_),
    .A2(_01755_),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08184_ (.A1(_01710_),
    .A2(_01756_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08185_ (.A1(_01700_),
    .A2(_01757_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08186_ (.A1(_01698_),
    .A2(_01758_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08187_ (.A1(_01695_),
    .A2(_01696_),
    .B(_01759_),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08188_ (.A1(_01695_),
    .A2(_01696_),
    .A3(_01759_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08189_ (.A1(_01761_),
    .A2(_01762_),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08190_ (.A1(_01693_),
    .A2(_01763_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08191_ (.A1(_00992_),
    .A2(_01764_),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08192_ (.A1(_01680_),
    .A2(_01682_),
    .B(_01691_),
    .C(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08193_ (.A1(_00138_),
    .A2(_01679_),
    .B(_01766_),
    .ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08194_ (.I(_00936_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08195_ (.A1(_01587_),
    .A2(_01589_),
    .B(_00779_),
    .C(_00788_),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08196_ (.A1(_01674_),
    .A2(_01768_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08197_ (.A1(_00930_),
    .A2(_00946_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08198_ (.A1(_01137_),
    .A2(_01769_),
    .B(_01771_),
    .ZN(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08199_ (.A1(_01767_),
    .A2(_01772_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08200_ (.A1(_01599_),
    .A2(_01659_),
    .A3(_01763_),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08201_ (.A1(_01695_),
    .A2(_01696_),
    .A3(_01759_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08202_ (.A1(_01692_),
    .A2(_01761_),
    .B(_01775_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08203_ (.A1(_01774_),
    .A2(_01776_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08204_ (.A1(_01700_),
    .A2(_01757_),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08205_ (.A1(_01698_),
    .A2(_01758_),
    .B(_01778_),
    .ZN(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08206_ (.A1(_00757_),
    .A2(_00775_),
    .A3(_01709_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08207_ (.A1(_01703_),
    .A2(_01708_),
    .B(_01780_),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08208_ (.A1(_01712_),
    .A2(_01755_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08209_ (.A1(_01710_),
    .A2(_01756_),
    .B(_01783_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08210_ (.A1(_01741_),
    .A2(_01753_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08211_ (.A1(_01741_),
    .A2(_01753_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08212_ (.A1(_01737_),
    .A2(_01785_),
    .B(_01786_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08213_ (.A1(_00789_),
    .A2(_01087_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08214_ (.A1(_01642_),
    .A2(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08215_ (.A1(_01742_),
    .A2(_01744_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08216_ (.A1(_01789_),
    .A2(_01790_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08217_ (.A1(_01787_),
    .A2(_01791_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08218_ (.A1(_00755_),
    .A2(_00931_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08219_ (.A1(_01793_),
    .A2(_01794_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08220_ (.A1(_01713_),
    .A2(_01734_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08221_ (.I(_01754_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08222_ (.A1(_01713_),
    .A2(_01734_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08223_ (.A1(_01796_),
    .A2(_01797_),
    .B(_01798_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08224_ (.A1(_01748_),
    .A2(_01752_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08225_ (.A1(_01748_),
    .A2(_01752_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08226_ (.A1(_01745_),
    .A2(_01800_),
    .B(_01801_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08227_ (.A1(_01728_),
    .A2(_01731_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08228_ (.A1(_01725_),
    .A2(_01732_),
    .B(_01804_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08229_ (.A1(net9),
    .A2(_00766_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08230_ (.A1(net8),
    .A2(_01223_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08231_ (.A1(_01788_),
    .A2(_01807_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08232_ (.A1(_01806_),
    .A2(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08233_ (.A1(_00903_),
    .A2(_00888_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08234_ (.A1(_01747_),
    .A2(_01751_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08235_ (.A1(_01648_),
    .A2(_01810_),
    .B1(_01811_),
    .B2(_01750_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08236_ (.A1(_00912_),
    .A2(_00875_),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08237_ (.A1(_01333_),
    .A2(_01096_),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08238_ (.A1(_01810_),
    .A2(_01813_),
    .A3(_01815_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08239_ (.A1(_01812_),
    .A2(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08240_ (.A1(_01809_),
    .A2(_01817_),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08241_ (.A1(_01802_),
    .A2(_01805_),
    .A3(_01818_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08242_ (.A1(_01721_),
    .A2(_01733_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08243_ (.A1(_01714_),
    .A2(_01720_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08244_ (.A1(_01048_),
    .A2(_00933_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08245_ (.A1(_00778_),
    .A2(_01161_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08246_ (.A1(net74),
    .A2(net16),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08247_ (.A1(_01714_),
    .A2(_01824_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08248_ (.A1(_01822_),
    .A2(_01823_),
    .B(_01826_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08249_ (.A1(_00913_),
    .A2(_01102_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08250_ (.A1(_00784_),
    .A2(net27),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08251_ (.A1(net71),
    .A2(_00828_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08252_ (.A1(_01829_),
    .A2(_01830_),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08253_ (.A1(_01828_),
    .A2(_01831_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08254_ (.A1(_01821_),
    .A2(_01827_),
    .A3(_01832_),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08255_ (.A1(_01723_),
    .A2(_01730_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08256_ (.A1(_00797_),
    .A2(_01156_),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08257_ (.A1(_01630_),
    .A2(_01835_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08258_ (.A1(_01729_),
    .A2(_01834_),
    .B(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08259_ (.A1(_01718_),
    .A2(_00845_),
    .B1(_00750_),
    .B2(_00785_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08260_ (.A1(_01552_),
    .A2(_01829_),
    .B1(_01839_),
    .B2(_01717_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08261_ (.A1(_00906_),
    .A2(_00892_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08262_ (.A1(_01259_),
    .A2(_01835_),
    .A3(_01841_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08263_ (.A1(_01840_),
    .A2(_01842_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08264_ (.A1(_01838_),
    .A2(_01843_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08265_ (.A1(_01833_),
    .A2(_01844_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08266_ (.A1(_01820_),
    .A2(_01845_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08267_ (.A1(_01819_),
    .A2(_01846_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08268_ (.A1(_01799_),
    .A2(_01848_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08269_ (.A1(_01795_),
    .A2(_01849_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08270_ (.A1(_01784_),
    .A2(_01850_),
    .Z(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08271_ (.A1(_01782_),
    .A2(_01851_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08272_ (.A1(_01779_),
    .A2(_01852_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08273_ (.A1(_01777_),
    .A2(_01853_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08274_ (.A1(_01767_),
    .A2(_01680_),
    .A3(_01688_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08275_ (.A1(_01680_),
    .A2(_01688_),
    .B(_01767_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08276_ (.A1(_05431_),
    .A2(_01856_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08277_ (.I(_00771_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08278_ (.A1(_00213_),
    .A2(_00934_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08279_ (.A1(_01767_),
    .A2(_01860_),
    .B(_05245_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08280_ (.A1(_01859_),
    .A2(_00130_),
    .B1(_00212_),
    .B2(_01666_),
    .C(_01861_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08281_ (.A1(_01685_),
    .A2(_00934_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08282_ (.A1(_00934_),
    .A2(_05280_),
    .B1(_01863_),
    .B2(_05282_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08283_ (.A1(_01685_),
    .A2(_04290_),
    .B(_01862_),
    .C(_01864_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08284_ (.A1(_01855_),
    .A2(_01857_),
    .B(_01865_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08285_ (.A1(_01345_),
    .A2(_01773_),
    .B1(_01854_),
    .B2(_01406_),
    .C(_01866_),
    .ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08286_ (.I(_00773_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08287_ (.A1(_01867_),
    .A2(_01863_),
    .A3(_01856_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08288_ (.A1(_01863_),
    .A2(_01856_),
    .B(_01867_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08289_ (.A1(_04097_),
    .A2(_01870_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08290_ (.I(_00940_),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08291_ (.A1(_00932_),
    .A2(_00935_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08292_ (.A1(_01873_),
    .A2(_01769_),
    .B(_00937_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08293_ (.A1(_01867_),
    .A2(_01874_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08294_ (.A1(_00939_),
    .A2(_00940_),
    .A3(_00938_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08295_ (.A1(_01867_),
    .A2(_00938_),
    .B(_01876_),
    .C(_01966_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08296_ (.A1(_01008_),
    .A2(_01875_),
    .B(_01877_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08297_ (.A1(_00939_),
    .A2(_01257_),
    .B1(_00584_),
    .B2(_01685_),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08298_ (.A1(_01859_),
    .A2(_01872_),
    .A3(_01193_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08299_ (.A1(_00418_),
    .A2(_00771_),
    .A3(_00940_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08300_ (.A1(_01859_),
    .A2(_01872_),
    .B(_04593_),
    .C(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08301_ (.A1(_01880_),
    .A2(_01881_),
    .A3(_01883_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08302_ (.A1(_01872_),
    .A2(_00421_),
    .B(_01878_),
    .C(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08303_ (.A1(_01779_),
    .A2(_01852_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08304_ (.A1(_01779_),
    .A2(_01852_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08305_ (.A1(_01777_),
    .A2(_01886_),
    .B(_01887_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08306_ (.A1(_01784_),
    .A2(_01850_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08307_ (.A1(_01782_),
    .A2(_01851_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08308_ (.A1(_00756_),
    .A2(_00931_),
    .A3(_01793_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08309_ (.A1(_01787_),
    .A2(_01791_),
    .B(_01892_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08310_ (.A1(_01799_),
    .A2(_01848_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08311_ (.A1(_01795_),
    .A2(_01849_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08312_ (.A1(_01894_),
    .A2(_01895_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08313_ (.A1(_01805_),
    .A2(_01818_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08314_ (.A1(_01805_),
    .A2(_01818_),
    .Z(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08315_ (.A1(_01802_),
    .A2(_01897_),
    .B(_01898_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08316_ (.A1(_01788_),
    .A2(_01807_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08317_ (.A1(_01806_),
    .A2(_01808_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08318_ (.A1(_01900_),
    .A2(_01902_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08319_ (.A1(_01899_),
    .A2(_01903_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08320_ (.A1(_00756_),
    .A2(_00770_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08321_ (.A1(_01904_),
    .A2(_01905_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08322_ (.A1(_01820_),
    .A2(_01845_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08323_ (.A1(_01819_),
    .A2(_01846_),
    .B(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08324_ (.A1(_01812_),
    .A2(_01816_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08325_ (.A1(_01809_),
    .A2(_01817_),
    .B(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08326_ (.A1(_01262_),
    .A2(_01835_),
    .A3(_01841_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08327_ (.A1(_01840_),
    .A2(_01911_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08328_ (.A1(_01838_),
    .A2(_01843_),
    .B(_01913_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08329_ (.A1(net10),
    .A2(_00766_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08330_ (.A1(net9),
    .A2(_00834_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08331_ (.A1(_01807_),
    .A2(_01916_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08332_ (.A1(_00780_),
    .A2(_00835_),
    .B1(_00850_),
    .B2(_00774_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08333_ (.A1(_01917_),
    .A2(_01918_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08334_ (.A1(_01915_),
    .A2(_01919_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08335_ (.A1(_01810_),
    .A2(_01815_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08336_ (.A1(_01334_),
    .A2(_00895_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08337_ (.A1(_01751_),
    .A2(_01922_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08338_ (.A1(_01813_),
    .A2(_01921_),
    .B(_01924_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08339_ (.A1(_00790_),
    .A2(_01071_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08340_ (.A1(_00918_),
    .A2(_00823_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08341_ (.A1(_01922_),
    .A2(_01927_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08342_ (.A1(_01926_),
    .A2(_01928_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08343_ (.A1(_01925_),
    .A2(_01929_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08344_ (.A1(_01925_),
    .A2(_01929_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08345_ (.A1(_01930_),
    .A2(_01931_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08346_ (.A1(_01920_),
    .A2(_01932_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08347_ (.A1(_01910_),
    .A2(_01914_),
    .A3(_01933_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08348_ (.A1(_01827_),
    .A2(_01832_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08349_ (.A1(_01827_),
    .A2(_01832_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08350_ (.A1(_01821_),
    .A2(_01935_),
    .A3(_01936_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08351_ (.A1(_01833_),
    .A2(_01844_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08352_ (.A1(_01937_),
    .A2(_01938_),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08353_ (.A1(net73),
    .A2(net27),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08354_ (.A1(net5),
    .A2(net75),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08355_ (.A1(_01824_),
    .A2(_01940_),
    .A3(_01941_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08356_ (.A1(_01826_),
    .A2(_01942_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08357_ (.A1(_00784_),
    .A2(_01030_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08358_ (.A1(net70),
    .A2(_01156_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08359_ (.A1(_01718_),
    .A2(_00870_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08360_ (.A1(_01945_),
    .A2(_01946_),
    .A3(_01947_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08361_ (.A1(_01943_),
    .A2(_01948_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08362_ (.A1(_01935_),
    .A2(_01949_),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08363_ (.A1(_00797_),
    .A2(_00892_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08364_ (.A1(_01835_),
    .A2(_01841_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08365_ (.A1(_01730_),
    .A2(_01951_),
    .B1(_01952_),
    .B2(_01261_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08366_ (.A1(_01719_),
    .A2(_01945_),
    .B1(_01831_),
    .B2(_01828_),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08367_ (.A1(_00904_),
    .A2(_00813_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08368_ (.A1(_00906_),
    .A2(_00809_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08369_ (.A1(_01951_),
    .A2(_01957_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08370_ (.A1(_01956_),
    .A2(_01958_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08371_ (.A1(_01954_),
    .A2(_01959_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08372_ (.A1(_01953_),
    .A2(_01960_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08373_ (.A1(_01950_),
    .A2(_01961_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08374_ (.A1(_01939_),
    .A2(_01962_),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08375_ (.A1(_01934_),
    .A2(_01963_),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08376_ (.A1(_01908_),
    .A2(_01964_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08377_ (.A1(_01906_),
    .A2(_01965_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08378_ (.A1(_01893_),
    .A2(_01896_),
    .A3(_01967_),
    .Z(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08379_ (.A1(_01889_),
    .A2(_01891_),
    .B(_01968_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08380_ (.A1(_01889_),
    .A2(_01891_),
    .A3(_01968_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08381_ (.A1(_01969_),
    .A2(_01970_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08382_ (.A1(_01888_),
    .A2(_01971_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08383_ (.A1(_00425_),
    .A2(_01972_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08384_ (.A1(_01869_),
    .A2(_01871_),
    .B(_01885_),
    .C(_01973_),
    .ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08385_ (.A1(_01899_),
    .A2(_01903_),
    .Z(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08386_ (.A1(_01904_),
    .A2(_01905_),
    .B(_01974_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08387_ (.A1(_01908_),
    .A2(_01964_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08388_ (.I(_01965_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08389_ (.A1(_01906_),
    .A2(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08390_ (.A1(_01977_),
    .A2(_01979_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08391_ (.A1(_01914_),
    .A2(_01933_),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08392_ (.A1(_01914_),
    .A2(_01933_),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08393_ (.A1(_01910_),
    .A2(_01981_),
    .B(_01982_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08394_ (.A1(_01915_),
    .A2(_01919_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08395_ (.A1(_01917_),
    .A2(_01984_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08396_ (.A1(_01983_),
    .A2(_01985_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08397_ (.A1(_01939_),
    .A2(_01962_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08398_ (.A1(_01934_),
    .A2(_01963_),
    .B(_01988_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08399_ (.A1(_01935_),
    .A2(_01949_),
    .Z(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08400_ (.A1(_01950_),
    .A2(_01961_),
    .B(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08401_ (.A1(_01826_),
    .A2(_01942_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08402_ (.A1(_01943_),
    .A2(_01948_),
    .B(_01992_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08403_ (.A1(_00772_),
    .A2(_00749_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08404_ (.A1(_01824_),
    .A2(_01941_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08405_ (.A1(_01822_),
    .A2(_01994_),
    .B1(_01995_),
    .B2(_01940_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08406_ (.A1(_00777_),
    .A2(_01030_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08407_ (.A1(_00933_),
    .A2(_01088_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08408_ (.A1(_01994_),
    .A2(_01997_),
    .A3(_01999_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08409_ (.A1(_01996_),
    .A2(_02000_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08410_ (.A1(_00914_),
    .A2(_00885_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08411_ (.A1(_00784_),
    .A2(_00870_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08412_ (.A1(_01718_),
    .A2(_00819_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08413_ (.A1(_02003_),
    .A2(_02004_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08414_ (.A1(_02002_),
    .A2(_02005_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08415_ (.A1(_02001_),
    .A2(_02006_),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08416_ (.A1(_01993_),
    .A2(_02007_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08417_ (.A1(_00798_),
    .A2(_00809_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08418_ (.A1(_01841_),
    .A2(_02010_),
    .B1(_01958_),
    .B2(_01956_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08419_ (.I(_02011_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08420_ (.A1(_01945_),
    .A2(_01947_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08421_ (.A1(_01830_),
    .A2(_02003_),
    .B1(_02013_),
    .B2(_01946_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08422_ (.A1(_01341_),
    .A2(_02010_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08423_ (.A1(_01334_),
    .A2(_00814_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08424_ (.A1(_02015_),
    .A2(_02016_),
    .Z(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08425_ (.A1(_02014_),
    .A2(_02017_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08426_ (.A1(_02012_),
    .A2(_02018_),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08427_ (.A1(_02008_),
    .A2(_02019_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08428_ (.A1(_01991_),
    .A2(_02021_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08429_ (.I(_02022_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08430_ (.A1(_01920_),
    .A2(_01932_),
    .B(_01930_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08431_ (.A1(_01954_),
    .A2(_01959_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08432_ (.A1(_01953_),
    .A2(_01960_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08433_ (.A1(_02025_),
    .A2(_02026_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08434_ (.A1(net11),
    .A2(_00767_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08435_ (.A1(net10),
    .A2(_00850_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08436_ (.A1(_01916_),
    .A2(_02029_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08437_ (.A1(_02028_),
    .A2(_02030_),
    .Z(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08438_ (.A1(_00918_),
    .A2(_00890_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08439_ (.A1(_01815_),
    .A2(_02033_),
    .B1(_01928_),
    .B2(_01926_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08440_ (.A1(_00780_),
    .A2(_01071_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08441_ (.A1(_00789_),
    .A2(_00824_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08442_ (.A1(_02033_),
    .A2(_02036_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08443_ (.A1(_02035_),
    .A2(_02037_),
    .Z(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08444_ (.A1(_02034_),
    .A2(_02038_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08445_ (.A1(_02032_),
    .A2(_02039_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08446_ (.A1(_02024_),
    .A2(_02027_),
    .A3(_02040_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08447_ (.A1(_02023_),
    .A2(_02041_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08448_ (.A1(_01989_),
    .A2(_02043_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08449_ (.A1(_01986_),
    .A2(_02044_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08450_ (.A1(_01975_),
    .A2(_01980_),
    .A3(_02045_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08451_ (.I(_01896_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08452_ (.A1(_02047_),
    .A2(_01967_),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08453_ (.A1(_02047_),
    .A2(_01967_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08454_ (.A1(_01893_),
    .A2(_02048_),
    .B(_02049_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08455_ (.A1(_02046_),
    .A2(_02050_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08456_ (.A1(_01889_),
    .A2(_01891_),
    .A3(_01968_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08457_ (.A1(_01887_),
    .A2(_01969_),
    .B(_02052_),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08458_ (.A1(_01776_),
    .A2(_02054_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08459_ (.A1(_01853_),
    .A2(_01969_),
    .A3(_01970_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08460_ (.A1(_01774_),
    .A2(_02055_),
    .B1(_02056_),
    .B2(_02054_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08461_ (.A1(_02051_),
    .A2(_02057_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08462_ (.I(_01872_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08463_ (.A1(_00939_),
    .A2(_02059_),
    .B(_01870_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08464_ (.A1(_01859_),
    .A2(_00585_),
    .B1(_02060_),
    .B2(_01028_),
    .C(_00588_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08465_ (.A1(_05115_),
    .A2(_02058_),
    .B(_02061_),
    .ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08466_ (.A1(_02046_),
    .A2(_02050_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08467_ (.A1(_01774_),
    .A2(_02055_),
    .B1(_02056_),
    .B2(_02054_),
    .C(_02051_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08468_ (.A1(_02062_),
    .A2(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08469_ (.A1(_01983_),
    .A2(_01985_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08470_ (.A1(_01989_),
    .A2(_02043_),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08471_ (.A1(_01986_),
    .A2(_02044_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08472_ (.A1(_02067_),
    .A2(_02068_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08473_ (.I(_02027_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08474_ (.A1(_02070_),
    .A2(_02040_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08475_ (.A1(_02070_),
    .A2(_02040_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08476_ (.A1(_02024_),
    .A2(_02071_),
    .B(_02072_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08477_ (.A1(_01916_),
    .A2(_02029_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08478_ (.A1(_02028_),
    .A2(_02030_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08479_ (.A1(_02075_),
    .A2(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08480_ (.A1(_02073_),
    .A2(_02077_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08481_ (.A1(_01991_),
    .A2(_02021_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08482_ (.A1(_02023_),
    .A2(_02041_),
    .B(_02079_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08483_ (.A1(_01993_),
    .A2(_02007_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08484_ (.A1(_02008_),
    .A2(_02019_),
    .B(_02081_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08485_ (.I(_01996_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08486_ (.A1(_02001_),
    .A2(_02006_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08487_ (.A1(_02083_),
    .A2(_02000_),
    .B(_02084_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08488_ (.A1(net75),
    .A2(_00844_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08489_ (.A1(_01994_),
    .A2(_01999_),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08490_ (.A1(_01824_),
    .A2(_02087_),
    .B1(_02088_),
    .B2(_01997_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08491_ (.A1(_00777_),
    .A2(_01102_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08492_ (.A1(net74),
    .A2(_00828_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08493_ (.A1(_02087_),
    .A2(_02091_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08494_ (.A1(_02090_),
    .A2(_02092_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08495_ (.A1(_02089_),
    .A2(_02093_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08496_ (.A1(_00785_),
    .A2(_00820_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08497_ (.A1(_00914_),
    .A2(_00811_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08498_ (.A1(_00793_),
    .A2(_00886_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08499_ (.A1(_02095_),
    .A2(_02097_),
    .A3(_02098_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08500_ (.A1(_02094_),
    .A2(_02099_),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08501_ (.I(_02100_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08502_ (.A1(_02086_),
    .A2(_02101_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08503_ (.I(_02102_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08504_ (.A1(_00799_),
    .A2(_00905_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08505_ (.A1(_01957_),
    .A2(_02104_),
    .B1(_02015_),
    .B2(_02016_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08506_ (.A1(_02003_),
    .A2(_02004_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08507_ (.A1(_02002_),
    .A2(_02005_),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08508_ (.A1(_02106_),
    .A2(_02108_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08509_ (.A1(_00919_),
    .A2(_00815_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08510_ (.A1(_01335_),
    .A2(_00806_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08511_ (.A1(_02104_),
    .A2(_02111_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08512_ (.A1(_02110_),
    .A2(_02112_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08513_ (.A1(_02109_),
    .A2(_02113_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08514_ (.A1(_02105_),
    .A2(_02114_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08515_ (.A1(_02103_),
    .A2(_02115_),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08516_ (.A1(_02082_),
    .A2(_02116_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08517_ (.A1(_02034_),
    .A2(_02038_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08518_ (.A1(_02032_),
    .A2(_02039_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08519_ (.A1(_02119_),
    .A2(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08520_ (.I(_02121_),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08521_ (.A1(_02014_),
    .A2(_02017_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08522_ (.A1(_02012_),
    .A2(_02018_),
    .B(_02123_),
    .ZN(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08523_ (.A1(net10),
    .A2(_00837_),
    .B1(_00852_),
    .B2(_00770_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08524_ (.A1(_00770_),
    .A2(_00837_),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08525_ (.A1(_02029_),
    .A2(_02126_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08526_ (.A1(_02125_),
    .A2(_02127_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08527_ (.A1(_00790_),
    .A2(_00890_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08528_ (.A1(_01927_),
    .A2(_02130_),
    .B1(_02037_),
    .B2(_02035_),
    .ZN(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08529_ (.A1(_00774_),
    .A2(_01072_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08530_ (.A1(_00781_),
    .A2(_00825_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08531_ (.A1(_02130_),
    .A2(_02133_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08532_ (.A1(_02132_),
    .A2(_02134_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08533_ (.A1(_02131_),
    .A2(_02135_),
    .Z(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08534_ (.A1(_02128_),
    .A2(_02136_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08535_ (.A1(_02122_),
    .A2(_02124_),
    .A3(_02137_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08536_ (.A1(_02117_),
    .A2(_02138_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08537_ (.A1(_02080_),
    .A2(_02139_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08538_ (.A1(_02078_),
    .A2(_02141_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08539_ (.A1(_02066_),
    .A2(_02069_),
    .A3(_02142_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08540_ (.A1(_01980_),
    .A2(_02045_),
    .Z(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08541_ (.A1(_01980_),
    .A2(_02045_),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08542_ (.A1(_01975_),
    .A2(_02144_),
    .B(_02145_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08543_ (.A1(_02143_),
    .A2(_02146_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08544_ (.A1(_02065_),
    .A2(_02147_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08545_ (.A1(_02065_),
    .A2(_02147_),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08546_ (.A1(_00671_),
    .A2(_02149_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08547_ (.A1(_02148_),
    .A2(_02150_),
    .B(_00674_),
    .ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08548_ (.I(_00951_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08549_ (.I(_02146_),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08550_ (.A1(_02143_),
    .A2(_02153_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08551_ (.A1(_02065_),
    .A2(_02147_),
    .B(_02154_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08552_ (.A1(_02067_),
    .A2(_02068_),
    .A3(_02142_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08553_ (.A1(_02067_),
    .A2(_02068_),
    .B(_02142_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08554_ (.A1(_02066_),
    .A2(_02156_),
    .B(_02157_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08555_ (.A1(_02080_),
    .A2(_02139_),
    .Z(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08556_ (.A1(_02078_),
    .A2(_02141_),
    .B(_02159_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08557_ (.I(_02114_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08558_ (.A1(_02105_),
    .A2(_02162_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08559_ (.A1(_02109_),
    .A2(_02113_),
    .B(_02163_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08560_ (.A1(_00781_),
    .A2(_00899_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08561_ (.A1(_02036_),
    .A2(_02165_),
    .B1(_02134_),
    .B2(_02132_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08562_ (.A1(_00931_),
    .A2(_01072_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08563_ (.A1(_02126_),
    .A2(_02165_),
    .A3(_02167_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08564_ (.A1(_02164_),
    .A2(_02166_),
    .A3(_02168_),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08565_ (.A1(_02073_),
    .A2(_02077_),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08566_ (.A1(_00920_),
    .A2(_00816_),
    .A3(_02112_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08567_ (.A1(_01271_),
    .A2(_02171_),
    .B(_01411_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08568_ (.A1(_01413_),
    .A2(_02171_),
    .B(_02173_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08569_ (.A1(_02170_),
    .A2(_02174_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08570_ (.I(_02082_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08571_ (.A1(_02176_),
    .A2(_02116_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08572_ (.A1(_02117_),
    .A2(_02138_),
    .B(_02177_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08573_ (.A1(_02124_),
    .A2(_02137_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08574_ (.A1(_02124_),
    .A2(_02137_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08575_ (.A1(_02122_),
    .A2(_02179_),
    .B(_02180_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08576_ (.A1(_00778_),
    .A2(_00822_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08577_ (.A1(_00933_),
    .A2(_00872_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08578_ (.A1(_00793_),
    .A2(_00811_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08579_ (.A1(_00772_),
    .A2(_00831_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08580_ (.A1(_01999_),
    .A2(_02186_),
    .B1(_02092_),
    .B2(_02090_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08581_ (.A1(_02184_),
    .A2(_02185_),
    .A3(_02187_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08582_ (.A1(_00786_),
    .A2(_00886_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08583_ (.A1(_02095_),
    .A2(_02098_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08584_ (.A1(_02004_),
    .A2(_02189_),
    .B1(_02190_),
    .B2(_02097_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08585_ (.A1(_00919_),
    .A2(_00807_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08586_ (.A1(_02189_),
    .A2(_02191_),
    .A3(_02192_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08587_ (.A1(_02182_),
    .A2(_02188_),
    .A3(_02193_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08588_ (.A1(_02086_),
    .A2(_02101_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08589_ (.A1(_02103_),
    .A2(_02115_),
    .B(_02196_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08590_ (.I(_02094_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08591_ (.A1(_02089_),
    .A2(_02093_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08592_ (.A1(_02198_),
    .A2(_02099_),
    .B(_02199_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08593_ (.A1(_00921_),
    .A2(_00905_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08594_ (.A1(_00790_),
    .A2(_00815_),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08595_ (.A1(_02186_),
    .A2(_02201_),
    .A3(_02202_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08596_ (.A1(_02197_),
    .A2(_02200_),
    .A3(_02203_),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08597_ (.A1(_02131_),
    .A2(_02135_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08598_ (.A1(_02128_),
    .A2(_02136_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08599_ (.A1(_02206_),
    .A2(_02207_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08600_ (.A1(_00775_),
    .A2(_00825_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08601_ (.A1(_02208_),
    .A2(_02209_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08602_ (.A1(_02195_),
    .A2(_02204_),
    .A3(_02210_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08603_ (.A1(_02127_),
    .A2(_02181_),
    .A3(_02211_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08604_ (.A1(_02175_),
    .A2(_02178_),
    .A3(_02212_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08605_ (.A1(_02169_),
    .A2(_02213_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08606_ (.A1(_02158_),
    .A2(_02160_),
    .A3(_02214_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08607_ (.A1(_02155_),
    .A2(_02215_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08608_ (.A1(_02155_),
    .A2(_02215_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08609_ (.A1(_02152_),
    .A2(_02217_),
    .A3(_02218_),
    .B(_00735_),
    .ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08610_ (.I(net47),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08611_ (.I(_02219_),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08612_ (.I(_02220_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08613_ (.I(_02221_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08614_ (.I(_02222_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08615_ (.I(_02223_),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08616_ (.I(net111),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08617_ (.I(_02225_),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08618_ (.I(_02227_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08619_ (.I(_02228_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08620_ (.I(_02229_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08621_ (.A1(_02222_),
    .A2(_02230_),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08622_ (.A1(_01498_),
    .A2(_02231_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08623_ (.I(net48),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08624_ (.I(_02233_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08625_ (.I(_02234_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08626_ (.I(_02235_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08627_ (.I(_02236_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08628_ (.I(_02230_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08629_ (.I(_02239_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08630_ (.A1(_02240_),
    .A2(_01890_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08631_ (.A1(_01825_),
    .A2(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _08632_ (.A1(_02238_),
    .A2(_01662_),
    .B1(_01738_),
    .B2(_02240_),
    .C1(_02224_),
    .C2(_02242_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08633_ (.A1(_02224_),
    .A2(_01249_),
    .B(_02232_),
    .C(_02243_),
    .ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08634_ (.I(_02220_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08635_ (.I(_02244_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08636_ (.A1(_02245_),
    .A2(_02240_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08637_ (.I(net112),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08638_ (.I(_02248_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08639_ (.I(_02249_),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08640_ (.I(_02250_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08641_ (.I(_02251_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08642_ (.A1(_02252_),
    .A2(_02235_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08643_ (.I(_02253_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08644_ (.I(net64),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08645_ (.A1(_02255_),
    .A2(net128),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08646_ (.I(_02256_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08647_ (.I(_02255_),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08648_ (.I(net128),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08649_ (.A1(_02259_),
    .A2(_02260_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08650_ (.A1(_02257_),
    .A2(_02261_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08651_ (.I(net127),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08652_ (.I(_02263_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08653_ (.I(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08654_ (.I(net63),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08655_ (.I(_02266_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08656_ (.I(_02267_),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08657_ (.I(_02268_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08658_ (.A1(_02265_),
    .A2(_02270_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08659_ (.I(net126),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08660_ (.I(_02272_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08661_ (.I(_02273_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08662_ (.I(net62),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08663_ (.A1(_02274_),
    .A2(_02275_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08664_ (.I(net123),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08665_ (.I(_02277_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08666_ (.I(net59),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08667_ (.I(_02279_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08668_ (.I(_02281_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08669_ (.I(_02282_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08670_ (.A1(_02278_),
    .A2(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08671_ (.I(net122),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08672_ (.I(_02285_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08673_ (.I(_02286_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08674_ (.I(_02287_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08675_ (.I(net58),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08676_ (.I(_02289_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08677_ (.I(_02290_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08678_ (.I(_02292_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08679_ (.A1(_02288_),
    .A2(_02293_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08680_ (.I(net121),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08681_ (.I(_02295_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08682_ (.I(_02296_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08683_ (.I(net57),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08684_ (.I(_02298_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08685_ (.I(_02299_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08686_ (.I(_02300_),
    .Z(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08687_ (.I(_02301_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08688_ (.A1(_02297_),
    .A2(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08689_ (.I(_02297_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08690_ (.I(_02301_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08691_ (.A1(_02305_),
    .A2(_02306_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08692_ (.I(net120),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08693_ (.I(_02308_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08694_ (.I(_02309_),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08695_ (.I(_02310_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08696_ (.I(net56),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08697_ (.I(_02312_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08698_ (.I(_02314_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08699_ (.I(_02315_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08700_ (.A1(_02311_),
    .A2(_02316_),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08701_ (.I(net119),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08702_ (.I(_02318_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08703_ (.I(_02319_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08704_ (.I(_02320_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08705_ (.I(net55),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08706_ (.I(_02322_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08707_ (.I(_02323_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08708_ (.I(_02325_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08709_ (.I(_02326_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08710_ (.I(_02327_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08711_ (.I(_02328_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08712_ (.A1(_02321_),
    .A2(_02329_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08713_ (.I(net118),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08714_ (.I(_02331_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08715_ (.I(_02332_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08716_ (.I(_02333_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08717_ (.I(_02334_),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08718_ (.I(_02336_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08719_ (.I(net54),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08720_ (.I(_02338_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08721_ (.I(_02339_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08722_ (.I(_02340_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08723_ (.I(_02341_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08724_ (.A1(_02337_),
    .A2(_02342_),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08725_ (.I(net117),
    .Z(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08726_ (.I(_02344_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08727_ (.I(_02345_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08728_ (.I(_02347_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08729_ (.I(_02348_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08730_ (.I(net53),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08731_ (.I(_02350_),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08732_ (.I(_02351_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08733_ (.I(_02352_),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08734_ (.A1(_02349_),
    .A2(_02353_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08735_ (.I(net116),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08736_ (.I(_02355_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08737_ (.I(_02356_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08738_ (.I(_02358_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08739_ (.I(_02359_),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08740_ (.I(net52),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08741_ (.I(_02361_),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08742_ (.I(_02362_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08743_ (.I(_02363_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08744_ (.A1(_02360_),
    .A2(_02364_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08745_ (.I(_02356_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08746_ (.A1(_02366_),
    .A2(_02363_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08747_ (.A1(_02365_),
    .A2(_02367_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08748_ (.I(net115),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08749_ (.I(_02370_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08750_ (.I(_02371_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08751_ (.I(net51),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08752_ (.I(_02373_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08753_ (.I(_02374_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08754_ (.I(_02375_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08755_ (.I(_02376_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08756_ (.A1(_02372_),
    .A2(_02377_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08757_ (.I(_02235_),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08758_ (.I(_02380_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08759_ (.A1(_02245_),
    .A2(_02239_),
    .B1(_02252_),
    .B2(_02381_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08760_ (.I(net114),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08761_ (.I(_02383_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08762_ (.I(net50),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08763_ (.I(_02385_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08764_ (.I(_02386_),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08765_ (.I(_02387_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08766_ (.I(_02388_),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08767_ (.A1(_02384_),
    .A2(_02389_),
    .B1(_02252_),
    .B2(_02381_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08768_ (.I(_02371_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08769_ (.I(_02392_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08770_ (.I(_02393_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08771_ (.A1(_02394_),
    .A2(_02376_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08772_ (.A1(_02394_),
    .A2(_02376_),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08773_ (.A1(_02395_),
    .A2(_02396_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08774_ (.A1(_02384_),
    .A2(_02389_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08775_ (.A1(_02382_),
    .A2(_02391_),
    .B(_02397_),
    .C(_02398_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08776_ (.A1(_02231_),
    .A2(_02253_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08777_ (.I(_02387_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08778_ (.A1(net114),
    .A2(_02402_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08779_ (.A1(_02400_),
    .A2(_02403_),
    .A3(_02397_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08780_ (.A1(_02378_),
    .A2(_02399_),
    .B(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08781_ (.I(_02348_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08782_ (.I(_02352_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08783_ (.A1(_02406_),
    .A2(_02407_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08784_ (.I(_02362_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08785_ (.A1(_02360_),
    .A2(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08786_ (.A1(_02369_),
    .A2(_02405_),
    .B(_02408_),
    .C(_02410_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08787_ (.I(_02342_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08788_ (.A1(_02337_),
    .A2(_02413_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08789_ (.A1(_02343_),
    .A2(_02354_),
    .A3(_02411_),
    .B(_02414_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08790_ (.A1(_02321_),
    .A2(_02329_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08791_ (.A1(_02311_),
    .A2(_02316_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08792_ (.A1(_02330_),
    .A2(_02415_),
    .B(_02416_),
    .C(_02417_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08793_ (.A1(_02307_),
    .A2(_02317_),
    .A3(_02418_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08794_ (.I(_02287_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08795_ (.A1(_02420_),
    .A2(_02292_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08796_ (.A1(_02420_),
    .A2(_02293_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08797_ (.A1(_02421_),
    .A2(_02422_),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08798_ (.A1(_02304_),
    .A2(_02419_),
    .A3(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08799_ (.A1(_02294_),
    .A2(_02425_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08800_ (.A1(_02278_),
    .A2(_02283_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08801_ (.A1(_02284_),
    .A2(_02426_),
    .B(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08802_ (.I(net125),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08803_ (.I(_02429_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08804_ (.I(_02430_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08805_ (.I(net61),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08806_ (.I(_02432_),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08807_ (.I(_02433_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08808_ (.A1(_02431_),
    .A2(_02435_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08809_ (.I(_02436_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08810_ (.I(_02435_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08811_ (.A1(_02431_),
    .A2(_02438_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08812_ (.A1(_02428_),
    .A2(_02437_),
    .B(_02439_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08813_ (.A1(_02274_),
    .A2(_02275_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08814_ (.A1(_02265_),
    .A2(_02268_),
    .B1(_02276_),
    .B2(_02440_),
    .C(_02441_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08815_ (.I(_02260_),
    .Z(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08816_ (.I(_02259_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08817_ (.I(_02444_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _08818_ (.A1(_02262_),
    .A2(_02271_),
    .A3(_02442_),
    .B1(_02443_),
    .B2(_02446_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08819_ (.A1(_02354_),
    .A2(_02408_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08820_ (.A1(_02369_),
    .A2(_02448_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08821_ (.A1(_02321_),
    .A2(_02328_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08822_ (.I(_02450_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08823_ (.I(_02340_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08824_ (.A1(_02336_),
    .A2(_02452_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08825_ (.A1(_02453_),
    .A2(_02414_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08826_ (.A1(_02404_),
    .A2(_02449_),
    .A3(_02451_),
    .A4(_02454_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08827_ (.A1(_02263_),
    .A2(_02268_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08828_ (.I(_02278_),
    .Z(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08829_ (.I(_02282_),
    .Z(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08830_ (.A1(_02458_),
    .A2(_02459_),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08831_ (.A1(_02304_),
    .A2(_02307_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08832_ (.I(net62),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08833_ (.I(_02462_),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08834_ (.A1(_02273_),
    .A2(_02463_),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08835_ (.A1(_02457_),
    .A2(_02460_),
    .A3(_02461_),
    .A4(_02464_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08836_ (.I(_02424_),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08837_ (.A1(_02257_),
    .A2(_02261_),
    .B(_02417_),
    .C(_02466_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08838_ (.A1(_02437_),
    .A2(_02468_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08839_ (.A1(_02455_),
    .A2(_02465_),
    .A3(_02469_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08840_ (.A1(_02447_),
    .A2(_02470_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08841_ (.I(_02471_),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08842_ (.A1(_02231_),
    .A2(_02472_),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08843_ (.A1(_02246_),
    .A2(_02254_),
    .A3(_02473_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08844_ (.I(_02252_),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08845_ (.I(_02248_),
    .Z(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08846_ (.I(net48),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08847_ (.A1(_02476_),
    .A2(_02477_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08848_ (.I(_02479_),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08849_ (.A1(_02475_),
    .A2(_02238_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08850_ (.A1(_04571_),
    .A2(_02480_),
    .B(_02481_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08851_ (.A1(_02222_),
    .A2(_02229_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08852_ (.I(_02248_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08853_ (.I(_02484_),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08854_ (.I(_02477_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08855_ (.I(_02486_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08856_ (.A1(_02485_),
    .A2(_02487_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08857_ (.I(_02488_),
    .Z(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08858_ (.A1(_02483_),
    .A2(_02490_),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08859_ (.A1(_02224_),
    .A2(_02475_),
    .B1(_02238_),
    .B2(_02240_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08860_ (.A1(_00951_),
    .A2(_02491_),
    .A3(_02492_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08861_ (.A1(_02475_),
    .A2(_00421_),
    .B1(_02482_),
    .B2(_04604_),
    .C(_02493_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08862_ (.I(_05375_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08863_ (.A1(_02483_),
    .A2(_02254_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08864_ (.A1(_02402_),
    .A2(_00233_),
    .B1(_00414_),
    .B2(_02381_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08865_ (.A1(_02224_),
    .A2(_00235_),
    .B1(_02480_),
    .B2(_00989_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08866_ (.A1(_02497_),
    .A2(_02498_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08867_ (.A1(_02495_),
    .A2(_02496_),
    .B(_02499_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08868_ (.A1(_04930_),
    .A2(_02474_),
    .B(_02494_),
    .C(_02501_),
    .ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08869_ (.I(_02383_),
    .Z(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08870_ (.I(_02502_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08871_ (.I(_02503_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08872_ (.I(_02504_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08873_ (.A1(_02223_),
    .A2(_02505_),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08874_ (.I(_02225_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08875_ (.I(_02507_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08876_ (.A1(_02508_),
    .A2(_02386_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08877_ (.A1(_02490_),
    .A2(_02491_),
    .A3(_02509_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08878_ (.I(net111),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08879_ (.I(_02512_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08880_ (.I(net50),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08881_ (.I(_02514_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08882_ (.A1(_02513_),
    .A2(_02515_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08883_ (.A1(_02483_),
    .A2(_02488_),
    .A3(_02516_),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08884_ (.I(_02516_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08885_ (.A1(_02480_),
    .A2(_02518_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08886_ (.A1(_02506_),
    .A2(_02511_),
    .A3(_02517_),
    .A4(_02519_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08887_ (.A1(_02511_),
    .A2(_02517_),
    .A3(_02519_),
    .B(_02506_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08888_ (.A1(_01113_),
    .A2(_02522_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08889_ (.I(_02502_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08890_ (.A1(_02524_),
    .A2(_02402_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08891_ (.A1(_02245_),
    .A2(_02239_),
    .B(_02254_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08892_ (.A1(_02475_),
    .A2(_02381_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08893_ (.A1(_02526_),
    .A2(_02527_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08894_ (.A1(_02525_),
    .A2(_02528_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08895_ (.A1(_02400_),
    .A2(_02472_),
    .A3(_02529_),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08896_ (.A1(_02400_),
    .A2(_02472_),
    .B(_02529_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08897_ (.A1(_05445_),
    .A2(_02531_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08898_ (.A1(_02530_),
    .A2(_02533_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08899_ (.A1(_02223_),
    .A2(_02239_),
    .A3(_02254_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08900_ (.A1(_02490_),
    .A2(_02535_),
    .B(_02525_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08901_ (.A1(_02490_),
    .A2(_02525_),
    .A3(_02535_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08902_ (.A1(_02536_),
    .A2(_02537_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08903_ (.I(_02504_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08904_ (.I(_02539_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08905_ (.A1(_02540_),
    .A2(_05497_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08906_ (.I(_02377_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08907_ (.A1(_02542_),
    .A2(_01338_),
    .B1(_02403_),
    .B2(_00238_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08908_ (.I(_02389_),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08909_ (.I(_01192_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08910_ (.A1(_02524_),
    .A2(_02545_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08911_ (.A1(_02545_),
    .A2(_01257_),
    .B1(_02546_),
    .B2(_02547_),
    .C1(_00968_),
    .C2(_02238_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08912_ (.A1(_02541_),
    .A2(_02544_),
    .A3(_02548_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08913_ (.A1(_02495_),
    .A2(_02538_),
    .B(_02549_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08914_ (.A1(_02520_),
    .A2(_02523_),
    .B(_02534_),
    .C(_02550_),
    .ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08915_ (.A1(_02382_),
    .A2(_02391_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08916_ (.A1(_02540_),
    .A2(_02545_),
    .B(_02551_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08917_ (.A1(_02525_),
    .A2(_02528_),
    .B(_02398_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08918_ (.I(_02470_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08919_ (.A1(_02447_),
    .A2(_02555_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08920_ (.I0(_02552_),
    .I1(_02554_),
    .S(_02556_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08921_ (.A1(_02397_),
    .A2(_02557_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08922_ (.A1(_02222_),
    .A2(_02394_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08923_ (.A1(_02375_),
    .A2(_02250_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08924_ (.I(_02560_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08925_ (.A1(_02479_),
    .A2(_02516_),
    .A3(_02561_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08926_ (.I(_02250_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08927_ (.A1(_02230_),
    .A2(_02376_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08928_ (.A1(_02388_),
    .A2(_02563_),
    .B(_02565_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08929_ (.A1(_02374_),
    .A2(_02249_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08930_ (.I(_02567_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08931_ (.A1(_02488_),
    .A2(_02518_),
    .A3(_02568_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08932_ (.A1(_02562_),
    .A2(_02566_),
    .A3(_02569_),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08933_ (.A1(_02517_),
    .A2(_02570_),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08934_ (.A1(_02559_),
    .A2(_02571_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08935_ (.A1(_02505_),
    .A2(_02236_),
    .A3(_02572_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08936_ (.A1(_02505_),
    .A2(_02236_),
    .B(_02572_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08937_ (.A1(_02573_),
    .A2(_02574_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08938_ (.A1(_02520_),
    .A2(_02576_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08939_ (.A1(_02547_),
    .A2(_02536_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08940_ (.A1(_02397_),
    .A2(_02578_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08941_ (.I(_05502_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08942_ (.I(_02364_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08943_ (.A1(_00395_),
    .A2(_02396_),
    .B(_02395_),
    .C(_00397_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08944_ (.A1(_02581_),
    .A2(_05191_),
    .B1(_05267_),
    .B2(_02402_),
    .C(_02582_),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08945_ (.I(_02394_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08946_ (.A1(_02584_),
    .A2(_00240_),
    .B1(_02396_),
    .B2(_01035_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08947_ (.A1(_02542_),
    .A2(_01238_),
    .B(_02583_),
    .C(_02585_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08948_ (.A1(_01152_),
    .A2(_02577_),
    .B1(_02579_),
    .B2(_02580_),
    .C(_02587_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08949_ (.A1(_00138_),
    .A2(_02558_),
    .B(_02588_),
    .ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08950_ (.A1(_02559_),
    .A2(_02571_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08951_ (.A1(_02223_),
    .A2(_02360_),
    .B1(_02584_),
    .B2(_02236_),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08952_ (.A1(_02359_),
    .A2(_02487_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08953_ (.I(_02591_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08954_ (.A1(_02559_),
    .A2(_02592_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08955_ (.A1(_02590_),
    .A2(_02593_),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08956_ (.I(_02225_),
    .Z(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08957_ (.A1(_02595_),
    .A2(_02361_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08958_ (.I(_02597_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08959_ (.A1(_02480_),
    .A2(_02518_),
    .A3(_02561_),
    .A4(_02598_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08960_ (.A1(_02230_),
    .A2(_02364_),
    .A3(_02388_),
    .A4(_02568_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08961_ (.A1(_02518_),
    .A2(_02561_),
    .B(_02598_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08962_ (.A1(_02562_),
    .A2(_02600_),
    .A3(_02601_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08963_ (.A1(_02517_),
    .A2(_02562_),
    .A3(_02566_),
    .A4(_02569_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08964_ (.A1(_02599_),
    .A2(_02602_),
    .B(_02603_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08965_ (.A1(_02603_),
    .A2(_02599_),
    .A3(_02602_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08966_ (.A1(_02604_),
    .A2(_02605_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08967_ (.A1(_02589_),
    .A2(_02594_),
    .A3(_02606_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08968_ (.A1(_02547_),
    .A2(_02608_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08969_ (.A1(_02520_),
    .A2(_02576_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08970_ (.A1(_02573_),
    .A2(_02610_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08971_ (.A1(_02609_),
    .A2(_02611_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08972_ (.I(_02369_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08973_ (.I(net51),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08974_ (.I(_02614_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08975_ (.A1(_02370_),
    .A2(_02615_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08976_ (.A1(_02584_),
    .A2(_02542_),
    .B1(_02547_),
    .B2(_02536_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08977_ (.A1(_02616_),
    .A2(_02617_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08978_ (.A1(_02613_),
    .A2(_02619_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08979_ (.I(_02353_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08980_ (.A1(_02581_),
    .A2(_00049_),
    .B1(_01368_),
    .B2(_02613_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08981_ (.A1(_02621_),
    .A2(_00983_),
    .B1(_02365_),
    .B2(_01265_),
    .C(_02622_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08982_ (.I(_02360_),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08983_ (.I(net52),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08984_ (.A1(_02355_),
    .A2(_02625_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08985_ (.I(_02626_),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08986_ (.A1(_02624_),
    .A2(_05280_),
    .B1(_05507_),
    .B2(_02542_),
    .C1(_02627_),
    .C2(_01577_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08987_ (.A1(_01118_),
    .A2(_02620_),
    .B(_02623_),
    .C(_02628_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08988_ (.I(_02404_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08989_ (.A1(_02631_),
    .A2(_02447_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08990_ (.A1(_02613_),
    .A2(_02405_),
    .A3(_02632_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08991_ (.A1(_04919_),
    .A2(_02633_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08992_ (.A1(_00425_),
    .A2(_02612_),
    .B(_02630_),
    .C(_02634_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08993_ (.I(_02635_),
    .ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08994_ (.A1(_02354_),
    .A2(_02408_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08995_ (.I(_02636_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08996_ (.A1(_02613_),
    .A2(_02405_),
    .B(_02410_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08997_ (.A1(_02624_),
    .A2(_02409_),
    .B(_02378_),
    .C(_02399_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08998_ (.A1(_02410_),
    .A2(_02640_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08999_ (.I(_02471_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09000_ (.I0(_02638_),
    .I1(_02641_),
    .S(_02642_),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09001_ (.A1(_02637_),
    .A2(_02643_),
    .B(_04756_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09002_ (.A1(_02637_),
    .A2(_02643_),
    .B(_02644_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09003_ (.A1(_02610_),
    .A2(_02609_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09004_ (.A1(_02573_),
    .A2(_02609_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09005_ (.A1(_02377_),
    .A2(_02383_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09006_ (.A1(_02593_),
    .A2(_02648_),
    .Z(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09007_ (.A1(_02603_),
    .A2(_02599_),
    .A3(_02602_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09008_ (.A1(_02594_),
    .A2(_02651_),
    .B(_02604_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09009_ (.A1(_02516_),
    .A2(_02567_),
    .A3(_02597_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09010_ (.A1(_02488_),
    .A2(_02509_),
    .A3(_02568_),
    .A4(_02597_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09011_ (.I(_02361_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09012_ (.I(net53),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09013_ (.I(_02656_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09014_ (.I(_02249_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09015_ (.A1(_02657_),
    .A2(_02658_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09016_ (.A1(_02507_),
    .A2(_02655_),
    .A3(_02568_),
    .A4(_02659_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09017_ (.I(_02660_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09018_ (.A1(_02227_),
    .A2(_02657_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09019_ (.A1(_02409_),
    .A2(_02563_),
    .B(_02663_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09020_ (.I(_02513_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09021_ (.A1(_02350_),
    .A2(_02484_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09022_ (.A1(_02665_),
    .A2(_02655_),
    .A3(_02560_),
    .A4(_02666_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09023_ (.A1(_02662_),
    .A2(_02664_),
    .A3(_02667_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09024_ (.A1(_02653_),
    .A2(_02654_),
    .A3(_02668_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09025_ (.A1(_02393_),
    .A2(_02387_),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09026_ (.I(_02219_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09027_ (.A1(_02671_),
    .A2(_02347_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09028_ (.A1(_02591_),
    .A2(_02673_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09029_ (.A1(_02670_),
    .A2(_02674_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09030_ (.A1(_02669_),
    .A2(_02675_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09031_ (.A1(_02649_),
    .A2(_02652_),
    .A3(_02676_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09032_ (.A1(_02590_),
    .A2(_02593_),
    .A3(_02604_),
    .A4(_02605_),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09033_ (.A1(_02590_),
    .A2(_02593_),
    .B1(_02604_),
    .B2(_02605_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09034_ (.A1(_02678_),
    .A2(_02679_),
    .B(_02589_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09035_ (.A1(_02589_),
    .A2(_02678_),
    .A3(_02679_),
    .ZN(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09036_ (.A1(_02524_),
    .A2(_02545_),
    .A3(_02680_),
    .B(_02681_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09037_ (.A1(_02677_),
    .A2(_02682_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09038_ (.A1(_02647_),
    .A2(_02684_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09039_ (.A1(_02646_),
    .A2(_02685_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09040_ (.A1(_01430_),
    .A2(_02686_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09041_ (.A1(_02616_),
    .A2(_02617_),
    .B(_02369_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09042_ (.A1(_02627_),
    .A2(_02688_),
    .B(_02636_),
    .ZN(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09043_ (.A1(_02627_),
    .A2(_02637_),
    .A3(_02688_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09044_ (.A1(_04485_),
    .A2(_02689_),
    .A3(_02690_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09045_ (.I(_01192_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09046_ (.A1(_02349_),
    .A2(_02407_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09047_ (.A1(_02413_),
    .A2(_04637_),
    .B1(_02692_),
    .B2(_02693_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09048_ (.A1(_02581_),
    .A2(_01410_),
    .B1(_02637_),
    .B2(_04593_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09049_ (.A1(_02621_),
    .A2(_05180_),
    .B(_02695_),
    .C(_02696_),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09050_ (.A1(_02406_),
    .A2(_00950_),
    .B(_02697_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09051_ (.A1(_02645_),
    .A2(_02687_),
    .A3(_02691_),
    .A4(_02698_),
    .ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09052_ (.I(_02471_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09053_ (.A1(_02406_),
    .A2(_02407_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09054_ (.A1(_02408_),
    .A2(_02410_),
    .A3(_02640_),
    .B(_02700_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09055_ (.A1(_02642_),
    .A2(_02701_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09056_ (.A1(_02354_),
    .A2(_02411_),
    .A3(_02699_),
    .B(_02702_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09057_ (.A1(_02454_),
    .A2(_02703_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09058_ (.A1(_02677_),
    .A2(_02682_),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09059_ (.A1(_02559_),
    .A2(_02592_),
    .A3(_02648_),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09060_ (.A1(_02652_),
    .A2(_02676_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09061_ (.A1(_02652_),
    .A2(_02676_),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09062_ (.A1(_02649_),
    .A2(_02708_),
    .B(_02709_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09063_ (.A1(_02592_),
    .A2(_02673_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09064_ (.A1(_02670_),
    .A2(_02674_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09065_ (.A1(_02711_),
    .A2(_02712_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09066_ (.A1(_02364_),
    .A2(_02383_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09067_ (.A1(_02713_),
    .A2(_02714_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09068_ (.A1(_02600_),
    .A2(_02601_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09069_ (.A1(_02653_),
    .A2(_02668_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09070_ (.A1(_02562_),
    .A2(_02717_),
    .A3(_02718_),
    .B1(_02669_),
    .B2(_02675_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09071_ (.A1(_02221_),
    .A2(_02334_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09072_ (.A1(_02345_),
    .A2(_02486_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09073_ (.I(_02514_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09074_ (.A1(_02358_),
    .A2(_02722_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09075_ (.A1(_02616_),
    .A2(_02721_),
    .A3(_02723_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09076_ (.A1(_02720_),
    .A2(_02724_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09077_ (.A1(_02653_),
    .A2(_02660_),
    .A3(_02664_),
    .A4(_02667_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09078_ (.A1(_02508_),
    .A2(_02452_),
    .A3(_02363_),
    .A4(_02666_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09079_ (.A1(_02228_),
    .A2(_02341_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09080_ (.A1(_02659_),
    .A2(_02729_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09081_ (.A1(_02508_),
    .A2(_02341_),
    .A3(_02409_),
    .A4(_02666_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09082_ (.A1(_02728_),
    .A2(_02730_),
    .A3(_02731_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09083_ (.A1(_02662_),
    .A2(_02727_),
    .A3(_02732_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09084_ (.A1(_02725_),
    .A2(_02733_),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09085_ (.A1(_02719_),
    .A2(_02734_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09086_ (.A1(_02716_),
    .A2(_02735_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09087_ (.A1(_02710_),
    .A2(_02736_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09088_ (.A1(_02707_),
    .A2(_02738_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09089_ (.A1(_02706_),
    .A2(_02739_),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09090_ (.A1(_02573_),
    .A2(_02609_),
    .A3(_02684_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09091_ (.A1(_02646_),
    .A2(_02685_),
    .B(_02741_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09092_ (.A1(_02740_),
    .A2(_02742_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09093_ (.I(_01727_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09094_ (.I(_02454_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09095_ (.A1(_02347_),
    .A2(_02351_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09096_ (.A1(_02745_),
    .A2(_02689_),
    .A3(_02746_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09097_ (.A1(_02689_),
    .A2(_02746_),
    .B(_02745_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09098_ (.A1(_02747_),
    .A2(_02749_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09099_ (.I(_04075_),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09100_ (.A1(net118),
    .A2(net54),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09101_ (.A1(_02621_),
    .A2(_01073_),
    .B1(_02752_),
    .B2(_01577_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09102_ (.I(_02328_),
    .Z(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09103_ (.A1(_02754_),
    .A2(_01417_),
    .B1(_05505_),
    .B2(_02452_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09104_ (.A1(_02413_),
    .A2(_05586_),
    .B1(_00133_),
    .B2(_02454_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09105_ (.A1(_02753_),
    .A2(_02755_),
    .A3(_02756_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09106_ (.A1(_02336_),
    .A2(_02744_),
    .B1(_02750_),
    .B2(_02751_),
    .C(_02757_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09107_ (.A1(_01345_),
    .A2(_02705_),
    .B1(_02743_),
    .B2(_01406_),
    .C(_02758_),
    .ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09108_ (.A1(_02414_),
    .A2(_02701_),
    .B(_02343_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09109_ (.A1(_02471_),
    .A2(_02760_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09110_ (.A1(_02415_),
    .A2(_02642_),
    .B(_02761_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09111_ (.A1(_02451_),
    .A2(_02762_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09112_ (.A1(_02706_),
    .A2(_02739_),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09113_ (.A1(_02740_),
    .A2(_02742_),
    .B(_02764_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09114_ (.A1(_02713_),
    .A2(_02714_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09115_ (.A1(_02719_),
    .A2(_02734_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09116_ (.A1(_02716_),
    .A2(_02735_),
    .B(_02767_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09117_ (.A1(_02345_),
    .A2(_02722_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09118_ (.A1(_02721_),
    .A2(_02723_),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09119_ (.A1(_02592_),
    .A2(_02770_),
    .B1(_02771_),
    .B2(_02616_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09120_ (.A1(_02352_),
    .A2(_02502_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09121_ (.A1(_02772_),
    .A2(_02773_),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09122_ (.A1(_02561_),
    .A2(_02598_),
    .A3(_02666_),
    .A4(_02729_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09123_ (.A1(_02662_),
    .A2(_02732_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09124_ (.A1(_02727_),
    .A2(_02775_),
    .A3(_02776_),
    .B1(_02733_),
    .B2(_02725_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09125_ (.A1(_02720_),
    .A2(_02724_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09126_ (.A1(_02221_),
    .A2(_02320_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09127_ (.A1(_02334_),
    .A2(_02235_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09128_ (.I(net119),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09129_ (.I(_02782_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09130_ (.A1(_02671_),
    .A2(_02783_),
    .A3(_02333_),
    .A4(_02234_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09131_ (.A1(_02779_),
    .A2(_02781_),
    .B(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09132_ (.A1(_02362_),
    .A2(_02370_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09133_ (.A1(_02366_),
    .A2(_02375_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09134_ (.A1(_02770_),
    .A2(_02786_),
    .A3(_02787_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09135_ (.A1(_02785_),
    .A2(_02788_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09136_ (.A1(_02778_),
    .A2(_02789_),
    .Z(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09137_ (.A1(_02598_),
    .A2(_02659_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09138_ (.I(_02512_),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09139_ (.I(_02248_),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09140_ (.A1(_02793_),
    .A2(_02339_),
    .A3(_02350_),
    .A4(_02794_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09141_ (.I(_02795_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09142_ (.A1(_02792_),
    .A2(_02796_),
    .Z(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09143_ (.A1(_02228_),
    .A2(_02325_),
    .B1(_02341_),
    .B2(_02485_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09144_ (.A1(_02595_),
    .A2(_02323_),
    .A3(_02340_),
    .A4(_02658_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09145_ (.A1(_02795_),
    .A2(_02799_),
    .Z(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09146_ (.A1(_02798_),
    .A2(_02800_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09147_ (.A1(_02797_),
    .A2(_02775_),
    .A3(_02801_),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09148_ (.A1(_02790_),
    .A2(_02803_),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09149_ (.A1(_02777_),
    .A2(_02804_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09150_ (.A1(_02774_),
    .A2(_02805_),
    .Z(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09151_ (.A1(_02766_),
    .A2(_02768_),
    .A3(_02806_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09152_ (.I(_02707_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09153_ (.A1(_02710_),
    .A2(_02736_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09154_ (.A1(_02808_),
    .A2(_02738_),
    .B(_02809_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09155_ (.A1(_02765_),
    .A2(_02807_),
    .A3(_02810_),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09156_ (.I(_05344_),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09157_ (.A1(_02451_),
    .A2(_02749_),
    .A3(_02752_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09158_ (.A1(_02749_),
    .A2(_02752_),
    .B(_02450_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09159_ (.A1(_02814_),
    .A2(_02815_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09160_ (.I(_02316_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09161_ (.A1(_02318_),
    .A2(_02322_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09162_ (.I(_02818_),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09163_ (.A1(_02754_),
    .A2(_04615_),
    .B1(_05591_),
    .B2(_02819_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09164_ (.A1(_02817_),
    .A2(_05589_),
    .B1(_05590_),
    .B2(_02413_),
    .C(_02820_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09165_ (.I(_05436_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09166_ (.A1(_02754_),
    .A2(_02822_),
    .B1(_05585_),
    .B2(_02451_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09167_ (.A1(_02821_),
    .A2(_02823_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09168_ (.A1(_02321_),
    .A2(_02744_),
    .B1(_02816_),
    .B2(_02751_),
    .C(_02825_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09169_ (.A1(_00137_),
    .A2(_02763_),
    .B1(_02811_),
    .B2(_02812_),
    .C(_02826_),
    .ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09170_ (.I(_02417_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09171_ (.A1(_02330_),
    .A2(_02415_),
    .B(_02416_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09172_ (.I(_02447_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09173_ (.A1(_02829_),
    .A2(_02455_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09174_ (.A1(_02827_),
    .A2(_02828_),
    .A3(_02830_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09175_ (.A1(_02807_),
    .A2(_02810_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09176_ (.A1(_02807_),
    .A2(_02810_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09177_ (.A1(_02765_),
    .A2(_02832_),
    .B(_02833_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09178_ (.A1(_02768_),
    .A2(_02806_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09179_ (.A1(_02768_),
    .A2(_02806_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09180_ (.A1(_02713_),
    .A2(_02714_),
    .A3(_02836_),
    .B(_02837_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09181_ (.A1(_02353_),
    .A2(_02539_),
    .A3(_02772_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09182_ (.A1(_02777_),
    .A2(_02804_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09183_ (.A1(_02774_),
    .A2(_02805_),
    .B(_02840_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09184_ (.A1(_02342_),
    .A2(_02384_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09185_ (.A1(_02778_),
    .A2(_02789_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09186_ (.A1(net117),
    .A2(_02373_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09187_ (.A1(_02770_),
    .A2(_02787_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09188_ (.A1(_02723_),
    .A2(_02844_),
    .B1(_02846_),
    .B2(_02786_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09189_ (.A1(_02843_),
    .A2(_02847_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09190_ (.A1(_02842_),
    .A2(_02848_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09191_ (.A1(_02730_),
    .A2(_02731_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09192_ (.A1(_02798_),
    .A2(_02800_),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09193_ (.A1(_02662_),
    .A2(_02797_),
    .A3(_02850_),
    .A4(_02851_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09194_ (.A1(_02790_),
    .A2(_02803_),
    .B(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09195_ (.A1(_02785_),
    .A2(_02788_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09196_ (.A1(_02656_),
    .A2(net115),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09197_ (.A1(_02626_),
    .A2(_02844_),
    .A3(_02855_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09198_ (.A1(_02782_),
    .A2(_02233_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09199_ (.A1(_02331_),
    .A2(_02385_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09200_ (.A1(_02220_),
    .A2(_02309_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09201_ (.A1(_02858_),
    .A2(_02859_),
    .A3(_02860_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09202_ (.A1(_02784_),
    .A2(_02857_),
    .A3(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09203_ (.A1(_02854_),
    .A2(_02862_),
    .Z(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09204_ (.I(_02799_),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09205_ (.I(_02864_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09206_ (.A1(_02796_),
    .A2(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09207_ (.A1(_02728_),
    .A2(_02798_),
    .A3(_02800_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09208_ (.A1(_02228_),
    .A2(_02314_),
    .A3(_02325_),
    .A4(_02485_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09209_ (.A1(_02229_),
    .A2(_02315_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09210_ (.A1(_02326_),
    .A2(_02251_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09211_ (.A1(_02864_),
    .A2(_02869_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09212_ (.A1(_02864_),
    .A2(_02869_),
    .B1(_02870_),
    .B2(_02871_),
    .C(_02872_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09213_ (.A1(_02866_),
    .A2(_02868_),
    .A3(_02873_),
    .Z(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09214_ (.A1(_02863_),
    .A2(_02874_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09215_ (.A1(_02853_),
    .A2(_02875_),
    .Z(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09216_ (.A1(_02849_),
    .A2(_02876_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09217_ (.A1(_02841_),
    .A2(_02877_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09218_ (.A1(_02839_),
    .A2(_02879_),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09219_ (.A1(_02838_),
    .A2(_02880_),
    .Z(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09220_ (.A1(_02835_),
    .A2(_02881_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09221_ (.A1(_02827_),
    .A2(_02815_),
    .A3(_02819_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09222_ (.A1(_02815_),
    .A2(_02819_),
    .B(_02827_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09223_ (.A1(_02883_),
    .A2(_02884_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09224_ (.A1(_00418_),
    .A2(_02311_),
    .B(_02827_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09225_ (.A1(_02817_),
    .A2(_01227_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09226_ (.A1(_02306_),
    .A2(_05435_),
    .B1(_02886_),
    .B2(_01123_),
    .C(_02887_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09227_ (.I(net120),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09228_ (.A1(_02890_),
    .A2(net56),
    .Z(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09229_ (.A1(_02310_),
    .A2(_00217_),
    .B1(_05332_),
    .B2(_02754_),
    .C1(_02891_),
    .C2(_05512_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09230_ (.A1(_02888_),
    .A2(_02892_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09231_ (.A1(_01152_),
    .A2(_02882_),
    .B1(_02885_),
    .B2(_02580_),
    .C(_02893_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09232_ (.A1(_00762_),
    .A2(_02831_),
    .B(_02894_),
    .ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09233_ (.A1(_02838_),
    .A2(_02880_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09234_ (.A1(_02835_),
    .A2(_02881_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09235_ (.A1(_02895_),
    .A2(_02896_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09236_ (.A1(_02841_),
    .A2(_02877_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09237_ (.A1(_02839_),
    .A2(_02879_),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09238_ (.A1(_02778_),
    .A2(_02789_),
    .A3(_02847_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09239_ (.A1(_02842_),
    .A2(_02848_),
    .B(_02901_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09240_ (.I(_02902_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09241_ (.A1(_02849_),
    .A2(_02876_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09242_ (.A1(_02853_),
    .A2(_02875_),
    .B(_02904_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09243_ (.A1(_02327_),
    .A2(_02503_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09244_ (.A1(_02854_),
    .A2(_02862_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09245_ (.A1(_02367_),
    .A2(_02844_),
    .Z(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09246_ (.A1(_02352_),
    .A2(_02584_),
    .A3(_02908_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09247_ (.A1(_02367_),
    .A2(_02844_),
    .B(_02909_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09248_ (.A1(_02907_),
    .A2(_02911_),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09249_ (.A1(_02906_),
    .A2(_02912_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09250_ (.A1(_02792_),
    .A2(_02796_),
    .A3(_02801_),
    .A4(_02873_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09251_ (.A1(_02863_),
    .A2(_02874_),
    .B(_02914_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09252_ (.A1(_02855_),
    .A2(_02908_),
    .Z(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09253_ (.A1(_02784_),
    .A2(_02861_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09254_ (.A1(_02784_),
    .A2(_02861_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09255_ (.A1(_02916_),
    .A2(_02917_),
    .B(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09256_ (.A1(_02347_),
    .A2(_02363_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09257_ (.A1(_02452_),
    .A2(_02372_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09258_ (.A1(_02351_),
    .A2(_02359_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09259_ (.A1(_02920_),
    .A2(_02922_),
    .A3(_02923_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09260_ (.A1(_02308_),
    .A2(_02233_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09261_ (.A1(_02671_),
    .A2(_02310_),
    .B1(_02320_),
    .B2(_02487_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09262_ (.A1(_02779_),
    .A2(_02925_),
    .B1(_02926_),
    .B2(_02859_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09263_ (.A1(_02332_),
    .A2(_02615_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09264_ (.A1(_02319_),
    .A2(_02722_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09265_ (.A1(_02925_),
    .A2(_02928_),
    .A3(_02929_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09266_ (.A1(_02927_),
    .A2(_02930_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09267_ (.A1(_02924_),
    .A2(_02931_),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09268_ (.A1(_02871_),
    .A2(_02870_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09269_ (.A1(_02796_),
    .A2(_02865_),
    .A3(_02869_),
    .A4(_02934_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09270_ (.A1(_02219_),
    .A2(net121),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09271_ (.I(_02312_),
    .Z(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09272_ (.I(_02476_),
    .Z(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09273_ (.A1(_02665_),
    .A2(_02937_),
    .A3(_02325_),
    .A4(_02938_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09274_ (.I(_02299_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09275_ (.A1(_02507_),
    .A2(_02940_),
    .A3(_02937_),
    .A4(_02938_),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09276_ (.A1(_02229_),
    .A2(_02301_),
    .B1(_02315_),
    .B2(_02251_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09277_ (.A1(_02939_),
    .A2(_02941_),
    .B(_02942_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09278_ (.A1(_02864_),
    .A2(_02869_),
    .A3(_02942_),
    .A4(_02941_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09279_ (.A1(_02939_),
    .A2(_02941_),
    .B1(_02944_),
    .B2(_02872_),
    .C(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09280_ (.A1(_02935_),
    .A2(_02936_),
    .A3(_02946_),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09281_ (.A1(_02919_),
    .A2(_02933_),
    .A3(_02947_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09282_ (.A1(_02915_),
    .A2(_02948_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09283_ (.A1(_02913_),
    .A2(_02949_),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09284_ (.A1(_02903_),
    .A2(_02905_),
    .A3(_02950_),
    .Z(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09285_ (.A1(_02898_),
    .A2(_02900_),
    .B(_02951_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09286_ (.A1(_02898_),
    .A2(_02900_),
    .A3(_02951_),
    .Z(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09287_ (.A1(_02952_),
    .A2(_02953_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09288_ (.A1(_02897_),
    .A2(_02955_),
    .Z(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09289_ (.I(_02461_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09290_ (.A1(_02891_),
    .A2(_02957_),
    .A3(_02884_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09291_ (.A1(_02891_),
    .A2(_02884_),
    .B(_02461_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09292_ (.A1(_02958_),
    .A2(_02959_),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09293_ (.A1(_02296_),
    .A2(_02300_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09294_ (.I(_02961_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09295_ (.A1(_02817_),
    .A2(_01410_),
    .B1(_02962_),
    .B2(_02692_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09296_ (.I(_02293_),
    .Z(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09297_ (.A1(_02964_),
    .A2(_05511_),
    .B1(_01418_),
    .B2(_02303_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09298_ (.A1(_02306_),
    .A2(_02822_),
    .B1(_05520_),
    .B2(_02957_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09299_ (.A1(_02963_),
    .A2(_02966_),
    .A3(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09300_ (.A1(_02297_),
    .A2(_01251_),
    .B1(_02960_),
    .B2(_01255_),
    .C(_02968_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09301_ (.A1(_02317_),
    .A2(_02418_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09302_ (.A1(_02311_),
    .A2(_02817_),
    .B1(_02330_),
    .B2(_02760_),
    .C(_02416_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09303_ (.A1(_02317_),
    .A2(_02971_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09304_ (.I0(_02970_),
    .I1(_02972_),
    .S(_02699_),
    .Z(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09305_ (.A1(_02957_),
    .A2(_02973_),
    .B(_01139_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09306_ (.A1(_02957_),
    .A2(_02973_),
    .B(_02974_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09307_ (.A1(_02812_),
    .A2(_02956_),
    .B(_02969_),
    .C(_02975_),
    .ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09308_ (.I(_05104_),
    .Z(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09309_ (.I(_02881_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09310_ (.A1(_02978_),
    .A2(_02955_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09311_ (.I(_02952_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09312_ (.A1(_02895_),
    .A2(_02980_),
    .B(_02953_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09313_ (.A1(_02835_),
    .A2(_02979_),
    .B(_02981_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09314_ (.A1(_02905_),
    .A2(_02950_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09315_ (.A1(_02905_),
    .A2(_02950_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09316_ (.A1(_02903_),
    .A2(_02983_),
    .B(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09317_ (.A1(_02328_),
    .A2(_02539_),
    .A3(_02912_),
    .Z(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09318_ (.A1(_02907_),
    .A2(_02911_),
    .B(_02987_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09319_ (.I(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09320_ (.A1(_02915_),
    .A2(_02948_),
    .Z(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09321_ (.A1(_02913_),
    .A2(_02949_),
    .B(_02990_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09322_ (.A1(_02316_),
    .A2(_02503_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09323_ (.A1(_02919_),
    .A2(_02933_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09324_ (.A1(_02920_),
    .A2(_02923_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09325_ (.A1(_02627_),
    .A2(_02693_),
    .B1(_02922_),
    .B2(_02994_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09326_ (.A1(_02993_),
    .A2(_02995_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09327_ (.A1(_02992_),
    .A2(_02996_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09328_ (.A1(_02919_),
    .A2(_02933_),
    .Z(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09329_ (.A1(_02936_),
    .A2(_02946_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09330_ (.A1(_02935_),
    .A2(_03000_),
    .Z(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09331_ (.A1(_02999_),
    .A2(_02947_),
    .B(_03001_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09332_ (.A1(_02927_),
    .A2(_02930_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09333_ (.A1(_02924_),
    .A2(_02931_),
    .B(_03003_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09334_ (.A1(_02308_),
    .A2(_02514_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09335_ (.I(_02308_),
    .Z(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09336_ (.A1(_02783_),
    .A2(_02386_),
    .B1(_02234_),
    .B2(_03006_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09337_ (.A1(_02858_),
    .A2(_03005_),
    .B1(_03007_),
    .B2(_02928_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09338_ (.A1(_02331_),
    .A2(_02625_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09339_ (.A1(_02318_),
    .A2(_02614_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09340_ (.A1(_03005_),
    .A2(_03010_),
    .A3(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09341_ (.A1(_03009_),
    .A2(_03012_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09342_ (.I(_02339_),
    .Z(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09343_ (.A1(_03014_),
    .A2(_02366_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09344_ (.A1(_02326_),
    .A2(_02392_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09345_ (.A1(_02746_),
    .A2(_03015_),
    .A3(_03016_),
    .Z(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09346_ (.A1(_03013_),
    .A2(_03017_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09347_ (.A1(_03004_),
    .A2(_03018_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09348_ (.A1(_02936_),
    .A2(_02946_),
    .B(_02945_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09349_ (.A1(_02244_),
    .A2(_02288_),
    .B1(_02305_),
    .B2(_02380_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09350_ (.A1(_02285_),
    .A2(net48),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09351_ (.I(_03023_),
    .Z(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09352_ (.A1(_02936_),
    .A2(_03024_),
    .Z(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09353_ (.A1(_03022_),
    .A2(_03025_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09354_ (.A1(_02507_),
    .A2(_02940_),
    .A3(_02937_),
    .A4(_02938_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09355_ (.A1(_02225_),
    .A2(_02289_),
    .A3(_02299_),
    .A4(_02476_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09356_ (.I(_03028_),
    .Z(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09357_ (.A1(_03027_),
    .A2(_03029_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09358_ (.A1(_02939_),
    .A2(_02941_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09359_ (.A1(_02665_),
    .A2(_02290_),
    .B1(_02300_),
    .B2(_02938_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09360_ (.A1(_03027_),
    .A2(_03029_),
    .B(_03033_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09361_ (.A1(_03032_),
    .A2(_03034_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09362_ (.A1(_03026_),
    .A2(_03031_),
    .A3(_03035_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09363_ (.A1(_03031_),
    .A2(_03035_),
    .B(_03026_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09364_ (.A1(_03036_),
    .A2(_03037_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09365_ (.A1(_03020_),
    .A2(_03021_),
    .A3(_03038_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09366_ (.A1(_03002_),
    .A2(_03039_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09367_ (.A1(_02991_),
    .A2(_02998_),
    .A3(_03040_),
    .Z(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09368_ (.A1(_02989_),
    .A2(_03042_),
    .Z(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09369_ (.A1(_02985_),
    .A2(_03043_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09370_ (.A1(_02985_),
    .A2(_03043_),
    .Z(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09371_ (.A1(_03044_),
    .A2(_03045_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09372_ (.A1(_02982_),
    .A2(_03046_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09373_ (.I(_02466_),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09374_ (.A1(_03048_),
    .A2(_02959_),
    .A3(_02961_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09375_ (.A1(_02959_),
    .A2(_02961_),
    .B(_02466_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09376_ (.A1(_01118_),
    .A2(_03050_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09377_ (.I(_02459_),
    .Z(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09378_ (.A1(_02964_),
    .A2(_04279_),
    .B1(_05321_),
    .B2(_03048_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09379_ (.A1(_03053_),
    .A2(_04334_),
    .B1(_02421_),
    .B2(_05320_),
    .C(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09380_ (.A1(_02420_),
    .A2(_02964_),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09381_ (.A1(_02420_),
    .A2(_01493_),
    .B1(_00968_),
    .B2(_02306_),
    .C1(_03056_),
    .C2(_02546_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09382_ (.A1(_03055_),
    .A2(_03057_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09383_ (.A1(_03049_),
    .A2(_03051_),
    .B(_03058_),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09384_ (.A1(_02304_),
    .A2(_02419_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09385_ (.A1(_02297_),
    .A2(_02303_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09386_ (.A1(_02304_),
    .A2(_02972_),
    .B(_03061_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09387_ (.I0(_03060_),
    .I1(_03062_),
    .S(_02699_),
    .Z(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09388_ (.A1(_03048_),
    .A2(_03064_),
    .B(_01139_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09389_ (.A1(_03048_),
    .A2(_03064_),
    .B(_03065_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09390_ (.A1(_02977_),
    .A2(_03047_),
    .B(_03059_),
    .C(_03066_),
    .ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09391_ (.I(_02460_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09392_ (.A1(_02288_),
    .A2(_02293_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09393_ (.A1(_02466_),
    .A2(_03062_),
    .B(_03068_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09394_ (.A1(_02642_),
    .A2(_03069_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09395_ (.A1(_02426_),
    .A2(_02699_),
    .B(_03070_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09396_ (.A1(_03067_),
    .A2(_03071_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09397_ (.A1(_02982_),
    .A2(_03046_),
    .B(_03044_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09398_ (.A1(_02998_),
    .A2(_03040_),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09399_ (.A1(_02991_),
    .A2(_03075_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09400_ (.A1(_02989_),
    .A2(_03042_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09401_ (.A1(_02993_),
    .A2(_02995_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09402_ (.A1(_02992_),
    .A2(_02996_),
    .B(_03078_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09403_ (.A1(_02999_),
    .A2(_02947_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09404_ (.A1(_03001_),
    .A2(_03080_),
    .B(_03039_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09405_ (.A1(_02998_),
    .A2(_03040_),
    .B(_03081_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09406_ (.A1(_02301_),
    .A2(_02503_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09407_ (.A1(_03004_),
    .A2(_03018_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09408_ (.A1(_02338_),
    .A2(_02344_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09409_ (.A1(_02746_),
    .A2(_03015_),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09410_ (.A1(_02923_),
    .A2(_03086_),
    .B1(_03016_),
    .B2(_03087_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09411_ (.A1(_03085_),
    .A2(_03088_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09412_ (.A1(_03083_),
    .A2(_03089_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09413_ (.A1(_03036_),
    .A2(_03037_),
    .B(_03021_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09414_ (.A1(_03021_),
    .A2(_03036_),
    .A3(_03037_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09415_ (.A1(_03020_),
    .A2(_03091_),
    .B(_03092_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09416_ (.A1(_03009_),
    .A2(_03012_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09417_ (.A1(_03013_),
    .A2(_03017_),
    .B(_03094_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09418_ (.A1(_02937_),
    .A2(_02371_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09419_ (.A1(_02322_),
    .A2(_02355_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09420_ (.A1(_03086_),
    .A2(_03098_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09421_ (.A1(_03097_),
    .A2(_03099_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09422_ (.A1(_02890_),
    .A2(_02614_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09423_ (.A1(_02319_),
    .A2(_02615_),
    .B1(_02515_),
    .B2(_02309_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09424_ (.A1(_02929_),
    .A2(_03101_),
    .B1(_03102_),
    .B2(_03010_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09425_ (.A1(net118),
    .A2(net53),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09426_ (.A1(_02318_),
    .A2(_02625_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09427_ (.A1(_03101_),
    .A2(_03104_),
    .A3(_03105_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09428_ (.A1(_03103_),
    .A2(_03107_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09429_ (.A1(_03100_),
    .A2(_03108_),
    .Z(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09430_ (.A1(_03096_),
    .A2(_03109_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09431_ (.A1(_03032_),
    .A2(_03034_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09432_ (.A1(_03026_),
    .A2(_03031_),
    .A3(_03035_),
    .B(_03111_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09433_ (.A1(net121),
    .A2(net50),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09434_ (.I(net123),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09435_ (.A1(_02219_),
    .A2(_03114_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09436_ (.A1(_03023_),
    .A2(_03113_),
    .A3(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09437_ (.A1(_03025_),
    .A2(_03116_),
    .Z(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09438_ (.I(net59),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09439_ (.I(_02289_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09440_ (.A1(_02595_),
    .A2(_03119_),
    .A3(_03120_),
    .A4(_02658_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09441_ (.A1(_03028_),
    .A2(_03121_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09442_ (.A1(_02665_),
    .A2(_02279_),
    .B1(_02290_),
    .B2(_02485_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09443_ (.A1(_02595_),
    .A2(_03120_),
    .A3(_02299_),
    .A4(_02484_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09444_ (.A1(_02512_),
    .A2(net59),
    .A3(net58),
    .A4(_02249_),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09445_ (.A1(_03124_),
    .A2(_03125_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09446_ (.A1(_03122_),
    .A2(_03123_),
    .A3(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09447_ (.A1(_03031_),
    .A2(_03118_),
    .A3(_03127_),
    .Z(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09448_ (.A1(_03112_),
    .A2(_03129_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09449_ (.A1(_03110_),
    .A2(_03130_),
    .Z(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09450_ (.A1(_03093_),
    .A2(_03131_),
    .Z(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09451_ (.A1(_03090_),
    .A2(_03132_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09452_ (.A1(_03079_),
    .A2(_03082_),
    .A3(_03133_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09453_ (.A1(_03076_),
    .A2(_03077_),
    .B(_03134_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09454_ (.A1(_03076_),
    .A2(_03077_),
    .A3(_03134_),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09455_ (.A1(_03135_),
    .A2(_03136_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09456_ (.A1(_03074_),
    .A2(_03137_),
    .B(_04442_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09457_ (.A1(_03074_),
    .A2(_03137_),
    .B(_03138_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09458_ (.A1(_03056_),
    .A2(_03067_),
    .A3(_03050_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09459_ (.A1(_03056_),
    .A2(_03050_),
    .B(_03067_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09460_ (.A1(_05375_),
    .A2(_03142_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09461_ (.A1(_03141_),
    .A2(_03143_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09462_ (.A1(_02964_),
    .A2(_00235_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09463_ (.A1(_02458_),
    .A2(_03053_),
    .A3(_00989_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09464_ (.I(_02438_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09465_ (.A1(_03147_),
    .A2(_00983_),
    .B1(_00234_),
    .B2(_02283_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09466_ (.A1(_03053_),
    .A2(_05437_),
    .B1(_01189_),
    .B2(_03067_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09467_ (.A1(_03145_),
    .A2(_03146_),
    .A3(_03148_),
    .A4(_03149_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09468_ (.A1(_02458_),
    .A2(_01251_),
    .B(_03144_),
    .C(_03151_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09469_ (.A1(_04930_),
    .A2(_03072_),
    .B(_03140_),
    .C(_03152_),
    .ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09470_ (.I(_03082_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09471_ (.A1(_03153_),
    .A2(_03133_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09472_ (.A1(_03153_),
    .A2(_03133_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09473_ (.A1(_03079_),
    .A2(_03154_),
    .B(_03155_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09474_ (.A1(_03004_),
    .A2(_03018_),
    .A3(_03088_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09475_ (.A1(_03083_),
    .A2(_03089_),
    .B(_03157_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09476_ (.I(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09477_ (.A1(_03093_),
    .A2(_03131_),
    .Z(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09478_ (.A1(_03090_),
    .A2(_03132_),
    .B(_03161_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09479_ (.A1(_02292_),
    .A2(_02502_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09480_ (.A1(_03096_),
    .A2(_03109_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09481_ (.A1(net55),
    .A2(net117),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09482_ (.A1(_03015_),
    .A2(_03165_),
    .B1(_03099_),
    .B2(_03097_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09483_ (.A1(_03164_),
    .A2(_03166_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09484_ (.A1(_03163_),
    .A2(_03167_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09485_ (.A1(_03112_),
    .A2(_03129_),
    .Z(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09486_ (.A1(_03110_),
    .A2(_03130_),
    .B(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09487_ (.A1(_03103_),
    .A2(_03107_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09488_ (.A1(_03100_),
    .A2(_03108_),
    .B(_03172_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09489_ (.A1(_03025_),
    .A2(_03116_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(net57),
    .A2(net115),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09491_ (.A1(net56),
    .A2(net116),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09492_ (.A1(_03165_),
    .A2(_03175_),
    .A3(_03176_),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09493_ (.A1(net120),
    .A2(net52),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09494_ (.A1(net119),
    .A2(net52),
    .B1(_02373_),
    .B2(net120),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09495_ (.A1(_03011_),
    .A2(_03178_),
    .B1(_03179_),
    .B2(_03104_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09496_ (.A1(net119),
    .A2(net53),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09497_ (.A1(_02752_),
    .A2(_03178_),
    .A3(_03181_),
    .Z(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09498_ (.A1(_03177_),
    .A2(_03180_),
    .A3(_03183_),
    .Z(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09499_ (.A1(_03174_),
    .A2(_03184_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09500_ (.A1(_03173_),
    .A2(_03185_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09501_ (.A1(_03122_),
    .A2(_03123_),
    .A3(_03126_),
    .B1(_03029_),
    .B2(_03027_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09502_ (.I(_03125_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09503_ (.A1(_03027_),
    .A2(_03029_),
    .A3(_03188_),
    .A4(_03123_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09504_ (.A1(_03118_),
    .A2(_03187_),
    .B(_03189_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09505_ (.A1(_03024_),
    .A2(_03115_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09506_ (.A1(_03024_),
    .A2(_03115_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09507_ (.A1(_03113_),
    .A2(_03191_),
    .B(_03192_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09508_ (.A1(_03114_),
    .A2(_02477_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09509_ (.A1(net121),
    .A2(_02614_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09510_ (.A1(_02286_),
    .A2(_02385_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09511_ (.A1(_03195_),
    .A2(_03196_),
    .A3(_03197_),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09512_ (.A1(_03194_),
    .A2(_03198_),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09513_ (.A1(_02244_),
    .A2(_02430_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09514_ (.A1(_02793_),
    .A2(net61),
    .A3(_03119_),
    .A4(_02484_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09515_ (.A1(_03188_),
    .A2(_03201_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09516_ (.A1(_02793_),
    .A2(net61),
    .A3(net59),
    .A4(_02794_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09517_ (.A1(_02227_),
    .A2(_02432_),
    .B1(_03119_),
    .B2(_02658_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09518_ (.A1(_03121_),
    .A2(_03203_),
    .B(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09519_ (.A1(_03202_),
    .A2(_03206_),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09520_ (.A1(_03126_),
    .A2(_03200_),
    .A3(_03207_),
    .Z(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09521_ (.A1(_03190_),
    .A2(_03199_),
    .A3(_03208_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09522_ (.A1(_03186_),
    .A2(_03209_),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09523_ (.A1(_03170_),
    .A2(_03210_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09524_ (.A1(_03168_),
    .A2(_03211_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09525_ (.A1(_03162_),
    .A2(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09526_ (.A1(_03159_),
    .A2(_03213_),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09527_ (.A1(_03159_),
    .A2(_03213_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09528_ (.A1(_03214_),
    .A2(_03216_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09529_ (.A1(_03156_),
    .A2(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09530_ (.I(_03136_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09531_ (.I(_03135_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09532_ (.A1(_03044_),
    .A2(_03220_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09533_ (.A1(_02835_),
    .A2(_02979_),
    .B1(_03219_),
    .B2(_03221_),
    .C(_02981_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09534_ (.A1(_03045_),
    .A2(_03135_),
    .B(_03219_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09535_ (.A1(_03222_),
    .A2(_03223_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09536_ (.A1(_03218_),
    .A2(_03224_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09537_ (.I(_02436_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09538_ (.A1(_02458_),
    .A2(_02459_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09539_ (.A1(_03227_),
    .A2(_03142_),
    .A3(_03228_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09540_ (.A1(_03142_),
    .A2(_03228_),
    .B(_02436_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09541_ (.A1(_01118_),
    .A2(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09542_ (.I(_02463_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09543_ (.A1(_00213_),
    .A2(_03147_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09544_ (.A1(_03227_),
    .A2(_03233_),
    .B(_04377_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09545_ (.A1(_03232_),
    .A2(_05589_),
    .B1(_05590_),
    .B2(_03053_),
    .C(_03234_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09546_ (.I(_02429_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09547_ (.I(_03236_),
    .Z(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09548_ (.A1(_03238_),
    .A2(_02438_),
    .Z(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09549_ (.A1(_03238_),
    .A2(_05583_),
    .B1(_03239_),
    .B2(_02546_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09550_ (.A1(_03147_),
    .A2(_00966_),
    .B(_03235_),
    .C(_03240_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09551_ (.A1(_03229_),
    .A2(_03231_),
    .B(_03241_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09552_ (.A1(_02284_),
    .A2(_03069_),
    .B(_02427_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09553_ (.A1(_02829_),
    .A2(_02555_),
    .B(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09554_ (.A1(_02428_),
    .A2(_02556_),
    .B(_03244_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09555_ (.A1(_03227_),
    .A2(_03245_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09556_ (.A1(_03227_),
    .A2(_03245_),
    .B(_03246_),
    .C(_01976_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09557_ (.A1(_02977_),
    .A2(_03225_),
    .B(_03242_),
    .C(_03247_),
    .ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09558_ (.I(_02464_),
    .Z(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09559_ (.A1(_02431_),
    .A2(_02438_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09560_ (.A1(_02436_),
    .A2(_03243_),
    .B(_03250_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09561_ (.A1(_02829_),
    .A2(_02555_),
    .B(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09562_ (.A1(_02440_),
    .A2(_02556_),
    .B(_03252_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09563_ (.I(_05444_),
    .Z(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09564_ (.A1(_03249_),
    .A2(_03253_),
    .B(_03254_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09565_ (.A1(_03249_),
    .A2(_03253_),
    .B(_03255_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09566_ (.A1(_03218_),
    .A2(_03222_),
    .A3(_03223_),
    .B1(_03217_),
    .B2(_03156_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09567_ (.A1(_03162_),
    .A2(_03212_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09568_ (.A1(_03096_),
    .A2(_03109_),
    .A3(_03166_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09569_ (.A1(_03163_),
    .A2(_03167_),
    .B(_03260_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09570_ (.I(_03170_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09571_ (.A1(_03262_),
    .A2(_03210_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09572_ (.A1(_03168_),
    .A2(_03211_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09573_ (.A1(_03263_),
    .A2(_03264_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09574_ (.A1(_02281_),
    .A2(_02384_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09575_ (.A1(_03174_),
    .A2(_03184_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09576_ (.A1(_03173_),
    .A2(_03185_),
    .B(_03267_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09577_ (.A1(net56),
    .A2(_02344_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09578_ (.A1(_03098_),
    .A2(_03270_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09579_ (.A1(_02327_),
    .A2(_02348_),
    .B(_03176_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09580_ (.A1(_03175_),
    .A2(_03271_),
    .A3(_03272_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09581_ (.A1(_03271_),
    .A2(_03273_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09582_ (.A1(_03268_),
    .A2(_03274_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09583_ (.A1(_03266_),
    .A2(_03275_),
    .Z(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09584_ (.I(_03190_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09585_ (.A1(_03199_),
    .A2(_03208_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09586_ (.A1(_03186_),
    .A2(_03209_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09587_ (.A1(_03277_),
    .A2(_03278_),
    .B(_03279_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09588_ (.A1(_03180_),
    .A2(_03183_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09589_ (.A1(_03180_),
    .A2(_03183_),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09590_ (.A1(_03177_),
    .A2(_03282_),
    .A3(_03283_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09591_ (.A1(_03282_),
    .A2(_03284_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09592_ (.A1(_03194_),
    .A2(_03198_),
    .Z(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09593_ (.I(_02289_),
    .Z(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09594_ (.A1(_03287_),
    .A2(_02370_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09595_ (.A1(_02298_),
    .A2(_02355_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09596_ (.A1(_03270_),
    .A2(_03289_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09597_ (.A1(_03288_),
    .A2(_03290_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09598_ (.A1(_02309_),
    .A2(_02657_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09599_ (.A1(_03178_),
    .A2(_03181_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09600_ (.A1(_02333_),
    .A2(_03014_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09601_ (.A1(_03105_),
    .A2(_03293_),
    .B1(_03294_),
    .B2(_03295_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09602_ (.A1(_02323_),
    .A2(_02332_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09603_ (.A1(_02319_),
    .A2(_02339_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09604_ (.A1(_03293_),
    .A2(_03297_),
    .A3(_03298_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09605_ (.A1(_03292_),
    .A2(_03296_),
    .A3(_03299_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09606_ (.A1(_03286_),
    .A2(_03300_),
    .Z(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09607_ (.A1(_03285_),
    .A2(_03301_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09608_ (.A1(_03200_),
    .A2(_03202_),
    .A3(_03206_),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09609_ (.A1(_03202_),
    .A2(_03206_),
    .B(_03200_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09610_ (.A1(_03124_),
    .A2(_03188_),
    .A3(_03304_),
    .A4(_03305_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09611_ (.A1(_03199_),
    .A2(_03208_),
    .B(_03306_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09612_ (.A1(net123),
    .A2(_02514_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09613_ (.A1(_02286_),
    .A2(_02722_),
    .B1(_02486_),
    .B2(_02277_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09614_ (.A1(_03024_),
    .A2(_03308_),
    .B1(_03309_),
    .B2(_03196_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09615_ (.I(_03310_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09616_ (.A1(_02295_),
    .A2(_02361_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09617_ (.A1(net122),
    .A2(_02373_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09618_ (.A1(_03308_),
    .A2(_03314_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09619_ (.A1(_03312_),
    .A2(_03315_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09620_ (.A1(_03311_),
    .A2(_03316_),
    .Z(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09621_ (.A1(_03188_),
    .A2(_03201_),
    .B(_03304_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09622_ (.A1(_02221_),
    .A2(_02273_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09623_ (.A1(_03236_),
    .A2(_02487_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09624_ (.A1(_02671_),
    .A2(_02272_),
    .A3(_03236_),
    .A4(_02234_),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09625_ (.A1(_03319_),
    .A2(_03320_),
    .B(_03321_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09626_ (.A1(_02508_),
    .A2(_02462_),
    .B1(_02433_),
    .B2(_02251_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09627_ (.I(_03323_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09628_ (.A1(_02227_),
    .A2(net62),
    .A3(_02432_),
    .A4(_02250_),
    .Z(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09629_ (.A1(_03201_),
    .A2(_03326_),
    .Z(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09630_ (.A1(_03322_),
    .A2(_03325_),
    .A3(_03327_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09631_ (.A1(_03325_),
    .A2(_03327_),
    .B(_03322_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09632_ (.A1(_03328_),
    .A2(_03329_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09633_ (.A1(_03317_),
    .A2(_03318_),
    .A3(_03330_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09634_ (.A1(_03307_),
    .A2(_03331_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09635_ (.A1(_03303_),
    .A2(_03332_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09636_ (.A1(_03276_),
    .A2(_03281_),
    .A3(_03333_),
    .Z(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09637_ (.I(_03334_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09638_ (.A1(_03265_),
    .A2(_03336_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09639_ (.A1(_03261_),
    .A2(_03337_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09640_ (.A1(_03259_),
    .A2(_03214_),
    .B(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09641_ (.A1(_03259_),
    .A2(_03214_),
    .A3(_03338_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09642_ (.A1(_03339_),
    .A2(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09643_ (.A1(_03257_),
    .A2(_03341_),
    .Z(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09644_ (.A1(_00244_),
    .A2(_03342_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09645_ (.A1(_03239_),
    .A2(_03230_),
    .B(_02464_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09646_ (.A1(_03239_),
    .A2(_03249_),
    .A3(_03230_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09647_ (.A1(_02751_),
    .A2(_03344_),
    .A3(_03345_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09648_ (.A1(_02274_),
    .A2(_01738_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09649_ (.A1(_02274_),
    .A2(_03232_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09650_ (.A1(_03147_),
    .A2(_04258_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09651_ (.I(_02270_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09652_ (.A1(_03351_),
    .A2(_00232_),
    .B1(_05384_),
    .B2(_02275_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09653_ (.A1(_05380_),
    .A2(_03349_),
    .B(_03350_),
    .C(_03352_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09654_ (.A1(_03232_),
    .A2(_00237_),
    .B1(_01189_),
    .B2(_03249_),
    .C(_03353_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09655_ (.A1(_03343_),
    .A2(_03347_),
    .A3(_03348_),
    .A4(_03354_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09656_ (.A1(_03256_),
    .A2(_03355_),
    .ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09657_ (.A1(_03218_),
    .A2(_03339_),
    .A3(_03340_),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09658_ (.A1(_03156_),
    .A2(_03217_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09659_ (.A1(_03358_),
    .A2(_03339_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09660_ (.A1(_03222_),
    .A2(_03223_),
    .A3(_03357_),
    .B1(_03359_),
    .B2(_03340_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09661_ (.A1(_02459_),
    .A2(_02540_),
    .A3(_03275_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09662_ (.A1(_03268_),
    .A2(_03274_),
    .B(_03361_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09663_ (.A1(_03281_),
    .A2(_03333_),
    .Z(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09664_ (.A1(_03281_),
    .A2(_03333_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09665_ (.A1(_03276_),
    .A2(_03363_),
    .B(_03364_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09666_ (.A1(_03286_),
    .A2(_03300_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09667_ (.A1(_03285_),
    .A2(_03301_),
    .B(_03366_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09668_ (.A1(_02303_),
    .A2(_02349_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09669_ (.A1(_03288_),
    .A2(_03290_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09670_ (.A1(_03176_),
    .A2(_03369_),
    .B(_03370_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09671_ (.A1(_03368_),
    .A2(_03371_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09672_ (.A1(_03368_),
    .A2(_03371_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09673_ (.A1(_03372_),
    .A2(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09674_ (.A1(_02435_),
    .A2(_02505_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09675_ (.A1(_03374_),
    .A2(_03375_),
    .Z(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09676_ (.I(_03307_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09677_ (.A1(_03377_),
    .A2(_03331_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09678_ (.A1(_03303_),
    .A2(_03332_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09679_ (.A1(_03379_),
    .A2(_03380_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09680_ (.A1(_03296_),
    .A2(_03299_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09681_ (.A1(_03296_),
    .A2(_03299_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09682_ (.A1(_03292_),
    .A2(_03382_),
    .B(_03383_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09683_ (.A1(_03311_),
    .A2(_03316_),
    .Z(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09684_ (.A1(_02281_),
    .A2(_02392_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09685_ (.I(_02344_),
    .Z(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09686_ (.A1(_03120_),
    .A2(_02940_),
    .A3(_03387_),
    .A4(_02358_),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09687_ (.A1(_02940_),
    .A2(_03387_),
    .B1(_02366_),
    .B2(_03287_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09688_ (.A1(_03388_),
    .A2(_03390_),
    .Z(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09689_ (.A1(_03386_),
    .A2(_03391_),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09690_ (.A1(_02890_),
    .A2(_02338_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09691_ (.A1(_02783_),
    .A2(_02340_),
    .B1(_02657_),
    .B2(_03006_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09692_ (.A1(_03181_),
    .A2(_03393_),
    .B1(_03394_),
    .B2(_03297_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09693_ (.A1(_02312_),
    .A2(_02332_),
    .Z(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09694_ (.A1(_02818_),
    .A2(_03393_),
    .A3(_03396_),
    .Z(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09695_ (.A1(_03395_),
    .A2(_03397_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09696_ (.A1(_03392_),
    .A2(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09697_ (.A1(_03385_),
    .A2(_03399_),
    .Z(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09698_ (.A1(_03384_),
    .A2(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09699_ (.A1(_03328_),
    .A2(_03329_),
    .B(_03318_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09700_ (.A1(_03318_),
    .A2(_03328_),
    .A3(_03329_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09701_ (.A1(_03317_),
    .A2(_03403_),
    .B(_03404_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09702_ (.A1(_02277_),
    .A2(_02615_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09703_ (.A1(_03197_),
    .A2(_03406_),
    .B1(_03315_),
    .B2(_03312_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09704_ (.A1(_02295_),
    .A2(_02350_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09705_ (.A1(_02286_),
    .A2(_02362_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09706_ (.A1(_03406_),
    .A2(_03408_),
    .A3(_03409_),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09707_ (.A1(_03321_),
    .A2(_03410_),
    .Z(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09708_ (.A1(_03407_),
    .A2(_03412_),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09709_ (.A1(_03201_),
    .A2(_03326_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09710_ (.A1(_03414_),
    .A2(_03328_),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09711_ (.A1(_02513_),
    .A2(_02266_),
    .A3(net62),
    .A4(_02794_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09712_ (.A1(_03326_),
    .A2(_03416_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09713_ (.A1(_02793_),
    .A2(_02266_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09714_ (.A1(_02275_),
    .A2(_02563_),
    .B(_03418_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09715_ (.A1(_03326_),
    .A2(_03416_),
    .Z(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09716_ (.A1(_03417_),
    .A2(_03419_),
    .A3(_03420_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09717_ (.A1(net126),
    .A2(_02233_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09718_ (.A1(_02429_),
    .A2(_02515_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09719_ (.A1(_02220_),
    .A2(_02263_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09720_ (.A1(_03423_),
    .A2(_03424_),
    .A3(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09721_ (.A1(_03421_),
    .A2(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09722_ (.A1(_03415_),
    .A2(_03427_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09723_ (.A1(_03405_),
    .A2(_03413_),
    .A3(_03428_),
    .Z(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09724_ (.A1(_03402_),
    .A2(_03429_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09725_ (.A1(_03381_),
    .A2(_03430_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09726_ (.A1(_03376_),
    .A2(_03431_),
    .Z(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09727_ (.A1(_03365_),
    .A2(_03432_),
    .Z(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09728_ (.A1(_03362_),
    .A2(_03434_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09729_ (.A1(_03265_),
    .A2(_03336_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09730_ (.A1(_03261_),
    .A2(_03337_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09731_ (.A1(_03436_),
    .A2(_03437_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09732_ (.A1(_03360_),
    .A2(_03435_),
    .A3(_03438_),
    .Z(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09733_ (.A1(_02265_),
    .A2(_02270_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09734_ (.A1(_03440_),
    .A2(_03344_),
    .A3(_03349_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09735_ (.A1(_03344_),
    .A2(_03349_),
    .B(_03440_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09736_ (.A1(_00964_),
    .A2(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09737_ (.A1(_00213_),
    .A2(_02270_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09738_ (.A1(_03440_),
    .A2(_03445_),
    .B(_05245_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09739_ (.A1(_02444_),
    .A2(_05589_),
    .B1(_00394_),
    .B2(_03232_),
    .C(_03446_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09740_ (.A1(_02264_),
    .A2(_03351_),
    .Z(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09741_ (.A1(_02264_),
    .A2(_05583_),
    .B1(_03448_),
    .B2(_02546_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09742_ (.A1(_03351_),
    .A2(_00966_),
    .B(_03447_),
    .C(_03449_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09743_ (.A1(_03441_),
    .A2(_03443_),
    .B(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09744_ (.A1(_02441_),
    .A2(_03251_),
    .B(_02276_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09745_ (.A1(_02276_),
    .A2(_02440_),
    .B(_02441_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09746_ (.A1(_03453_),
    .A2(_02829_),
    .A3(_02555_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09747_ (.A1(_02556_),
    .A2(_03452_),
    .B(_03454_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09748_ (.A1(_02457_),
    .A2(_03456_),
    .B(_01139_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09749_ (.A1(_02457_),
    .A2(_03456_),
    .B(_03457_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09750_ (.A1(_02977_),
    .A2(_03439_),
    .B(_03451_),
    .C(_03458_),
    .ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09751_ (.A1(_02446_),
    .A2(_02443_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09752_ (.A1(_02271_),
    .A2(_02442_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09753_ (.A1(_03440_),
    .A2(_03452_),
    .B(_02271_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09754_ (.A1(_02262_),
    .A2(_03461_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09755_ (.A1(_03459_),
    .A2(_03460_),
    .B1(_02472_),
    .B2(_03462_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09756_ (.A1(_04919_),
    .A2(_03463_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09757_ (.A1(_02446_),
    .A2(_00414_),
    .B1(_04215_),
    .B2(_02257_),
    .C1(_00235_),
    .C2(_03351_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09758_ (.A1(_04571_),
    .A2(_02257_),
    .B(_02261_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09759_ (.A1(_02443_),
    .A2(_00988_),
    .B1(_03467_),
    .B2(_00238_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09760_ (.A1(_03466_),
    .A2(_03468_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09761_ (.A1(_03464_),
    .A2(_03469_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09762_ (.A1(_03374_),
    .A2(_03375_),
    .B(_03373_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09763_ (.A1(_03379_),
    .A2(_03380_),
    .B(_03430_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09764_ (.A1(_03376_),
    .A2(_03431_),
    .B(_03472_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09765_ (.A1(_03385_),
    .A2(_03399_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09766_ (.A1(_03384_),
    .A2(_03401_),
    .B(_03474_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09767_ (.A1(_03386_),
    .A2(_03391_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09768_ (.A1(_03388_),
    .A2(_03477_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09769_ (.A1(_03475_),
    .A2(_03478_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09770_ (.A1(_03475_),
    .A2(_03478_),
    .Z(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09771_ (.A1(_03479_),
    .A2(_03480_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09772_ (.A1(_02463_),
    .A2(_02504_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09773_ (.A1(_03481_),
    .A2(_03482_),
    .Z(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09774_ (.A1(_03413_),
    .A2(_03428_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09775_ (.A1(_03413_),
    .A2(_03428_),
    .Z(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09776_ (.A1(_03405_),
    .A2(_03484_),
    .A3(_03485_),
    .B1(_03429_),
    .B2(_03402_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09777_ (.A1(_03395_),
    .A2(_03397_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09778_ (.A1(_03392_),
    .A2(_03398_),
    .B(_03488_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09779_ (.I(_03412_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09780_ (.A1(_02245_),
    .A2(_02431_),
    .A3(_03423_),
    .A4(_03410_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09781_ (.A1(_03407_),
    .A2(_03490_),
    .B(_03491_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09782_ (.A1(_02433_),
    .A2(_02371_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09783_ (.A1(_03119_),
    .A2(_03120_),
    .A3(_02345_),
    .A4(_02356_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09784_ (.A1(_03287_),
    .A2(_03387_),
    .B1(_02358_),
    .B2(_02279_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09785_ (.A1(_03494_),
    .A2(_03495_),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09786_ (.A1(_03493_),
    .A2(_03496_),
    .Z(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09787_ (.A1(_02818_),
    .A2(_03393_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09788_ (.A1(_02890_),
    .A2(_02322_),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09789_ (.A1(_03298_),
    .A2(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09790_ (.A1(_03499_),
    .A2(_03396_),
    .B(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09791_ (.A1(_02298_),
    .A2(_02331_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09792_ (.A1(_02312_),
    .A2(_02782_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09793_ (.A1(_03500_),
    .A2(_03503_),
    .A3(_03504_),
    .Z(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09794_ (.A1(_03502_),
    .A2(_03505_),
    .Z(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09795_ (.A1(_03497_),
    .A2(_03506_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09796_ (.A1(_03492_),
    .A2(_03507_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09797_ (.A1(_03489_),
    .A2(_03508_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09798_ (.A1(_03415_),
    .A2(_03427_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09799_ (.A1(_03413_),
    .A2(_03428_),
    .B(_03511_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09800_ (.A1(_03417_),
    .A2(_03419_),
    .A3(_03420_),
    .A4(_03426_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09801_ (.A1(_03417_),
    .A2(_03513_),
    .Z(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09802_ (.A1(net63),
    .A2(net112),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09803_ (.A1(net47),
    .A2(net128),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09804_ (.A1(_02512_),
    .A2(net64),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09805_ (.A1(_03515_),
    .A2(_03516_),
    .A3(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09806_ (.A1(_03416_),
    .A2(_03518_),
    .Z(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09807_ (.A1(net127),
    .A2(_02477_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09808_ (.A1(net125),
    .A2(_02374_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09809_ (.A1(_02272_),
    .A2(_02515_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09810_ (.A1(_03521_),
    .A2(_03522_),
    .A3(_03523_),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09811_ (.A1(_03519_),
    .A2(_03524_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09812_ (.A1(_03514_),
    .A2(_03525_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09813_ (.A1(_03114_),
    .A2(_02625_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09814_ (.A1(_03406_),
    .A2(_03409_),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09815_ (.A1(_03314_),
    .A2(_03527_),
    .B1(_03528_),
    .B2(_03408_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09816_ (.A1(_03423_),
    .A2(_03425_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09817_ (.A1(_03319_),
    .A2(_03521_),
    .B1(_03530_),
    .B2(_03424_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09818_ (.A1(_02296_),
    .A2(_03014_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09819_ (.A1(_02285_),
    .A2(_02656_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09820_ (.A1(_03527_),
    .A2(_03534_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09821_ (.A1(_03533_),
    .A2(_03535_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09822_ (.A1(_03532_),
    .A2(_03536_),
    .Z(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09823_ (.A1(_03529_),
    .A2(_03537_),
    .Z(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09824_ (.A1(_03526_),
    .A2(_03538_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09825_ (.A1(_03512_),
    .A2(_03539_),
    .Z(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09826_ (.A1(_03510_),
    .A2(_03540_),
    .Z(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09827_ (.A1(_03486_),
    .A2(_03541_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09828_ (.A1(_03483_),
    .A2(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09829_ (.A1(_03473_),
    .A2(_03544_),
    .Z(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09830_ (.A1(_03471_),
    .A2(_03545_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09831_ (.I(_03546_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09832_ (.A1(_03365_),
    .A2(_03432_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09833_ (.A1(_03362_),
    .A2(_03434_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09834_ (.A1(_03548_),
    .A2(_03549_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09835_ (.A1(_03547_),
    .A2(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09836_ (.A1(_03547_),
    .A2(_03550_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09837_ (.I(_03552_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09838_ (.A1(_03551_),
    .A2(_03554_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09839_ (.A1(_03436_),
    .A2(_03437_),
    .A3(_03435_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09840_ (.A1(_03436_),
    .A2(_03437_),
    .B(_03435_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09841_ (.A1(_03360_),
    .A2(_03556_),
    .B(_03557_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09842_ (.A1(_03555_),
    .A2(_03558_),
    .Z(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09843_ (.A1(_03448_),
    .A2(_03442_),
    .B(_02262_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09844_ (.A1(_02262_),
    .A2(_03448_),
    .A3(_03442_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09845_ (.A1(_00979_),
    .A2(_03561_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09846_ (.A1(_00425_),
    .A2(_03559_),
    .B1(_03560_),
    .B2(_03562_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09847_ (.A1(_03470_),
    .A2(_03563_),
    .ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09848_ (.A1(_03481_),
    .A2(_03482_),
    .B(_03480_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09849_ (.A1(_03486_),
    .A2(_03541_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09850_ (.A1(_03483_),
    .A2(_03543_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09851_ (.A1(_03566_),
    .A2(_03567_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09852_ (.A1(_03512_),
    .A2(_03539_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09853_ (.A1(_03510_),
    .A2(_03540_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09854_ (.A1(_03569_),
    .A2(_03570_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09855_ (.A1(_03514_),
    .A2(_03525_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09856_ (.A1(_03526_),
    .A2(_03538_),
    .B(_03572_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09857_ (.I(_03416_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09858_ (.A1(_03575_),
    .A2(_03518_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09859_ (.A1(_03519_),
    .A2(_03524_),
    .B(_03576_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09860_ (.A1(_02255_),
    .A2(_02476_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09861_ (.A1(net128),
    .A2(_02486_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09862_ (.A1(_02479_),
    .A2(_02256_),
    .B1(_03578_),
    .B2(_03579_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09863_ (.A1(_02513_),
    .A2(_02255_),
    .B1(_02266_),
    .B2(_02794_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09864_ (.A1(_03418_),
    .A2(_03578_),
    .B1(_03581_),
    .B2(_03516_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09865_ (.A1(_03580_),
    .A2(_03582_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09866_ (.A1(net127),
    .A2(_02385_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09867_ (.A1(net126),
    .A2(_02374_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09868_ (.A1(_03584_),
    .A2(_03586_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09869_ (.A1(_02429_),
    .A2(_02655_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09870_ (.A1(_03587_),
    .A2(_03588_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09871_ (.A1(_03583_),
    .A2(_03589_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09872_ (.A1(_03577_),
    .A2(_03590_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09873_ (.A1(_03114_),
    .A2(_02656_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09874_ (.A1(_03409_),
    .A2(_03592_),
    .B1(_03535_),
    .B2(_03533_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09875_ (.I(_03593_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09876_ (.A1(_03521_),
    .A2(_03523_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09877_ (.A1(_03423_),
    .A2(_03584_),
    .B1(_03595_),
    .B2(_03522_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09878_ (.A1(_02295_),
    .A2(_02323_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09879_ (.A1(_02285_),
    .A2(_02338_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09880_ (.A1(_03592_),
    .A2(_03599_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09881_ (.A1(_03598_),
    .A2(_03600_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09882_ (.A1(_03597_),
    .A2(_03601_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09883_ (.A1(_03594_),
    .A2(_03602_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09884_ (.A1(_03591_),
    .A2(_03603_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09885_ (.A1(_03573_),
    .A2(_03604_),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09886_ (.A1(_03497_),
    .A2(_03506_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09887_ (.A1(_03502_),
    .A2(_03505_),
    .B(_03606_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09888_ (.I(_03529_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09889_ (.I(_03536_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09890_ (.A1(_03532_),
    .A2(_03610_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09891_ (.A1(_03609_),
    .A2(_03537_),
    .B(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09892_ (.A1(_02462_),
    .A2(_02392_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09893_ (.A1(_02279_),
    .A2(_03387_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09894_ (.A1(_02432_),
    .A2(_02356_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09895_ (.A1(_03614_),
    .A2(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09896_ (.A1(_03613_),
    .A2(_03616_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09897_ (.A1(_03006_),
    .A2(_02314_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09898_ (.A1(_03500_),
    .A2(_03504_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09899_ (.A1(_03619_),
    .A2(_02819_),
    .B1(_03503_),
    .B2(_03620_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09900_ (.A1(_02298_),
    .A2(_02782_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09901_ (.A1(_02891_),
    .A2(_03622_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09902_ (.A1(_03287_),
    .A2(_02333_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09903_ (.A1(_03623_),
    .A2(_03624_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09904_ (.A1(_03621_),
    .A2(_03625_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09905_ (.I(_03626_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09906_ (.A1(_03617_),
    .A2(_03627_),
    .Z(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09907_ (.A1(_03612_),
    .A2(_03628_),
    .Z(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09908_ (.A1(_03608_),
    .A2(_03630_),
    .Z(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09909_ (.A1(_03605_),
    .A2(_03631_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09910_ (.A1(_03571_),
    .A2(_03632_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09911_ (.I(_03508_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09912_ (.A1(_03492_),
    .A2(_03507_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09913_ (.A1(_03489_),
    .A2(_03634_),
    .B(_03635_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09914_ (.A1(_03493_),
    .A2(_03496_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09915_ (.A1(_03494_),
    .A2(_03637_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09916_ (.A1(_03636_),
    .A2(_03638_),
    .Z(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09917_ (.A1(_02267_),
    .A2(_02504_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09918_ (.A1(_03639_),
    .A2(_03641_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09919_ (.A1(_03633_),
    .A2(_03642_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09920_ (.A1(_03568_),
    .A2(_03643_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09921_ (.A1(_03565_),
    .A2(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09922_ (.A1(_03473_),
    .A2(_03544_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09923_ (.A1(_03471_),
    .A2(_03545_),
    .B(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09924_ (.A1(_03645_),
    .A2(_03647_),
    .Z(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09925_ (.A1(_03552_),
    .A2(_03558_),
    .B(_03551_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09926_ (.A1(_03648_),
    .A2(_03649_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09927_ (.A1(_03648_),
    .A2(_03649_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09928_ (.A1(_00671_),
    .A2(_03652_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09929_ (.A1(_02444_),
    .A2(_02443_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09930_ (.A1(_03654_),
    .A2(_03560_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09931_ (.A1(_02444_),
    .A2(_00585_),
    .B1(_03655_),
    .B2(_02580_),
    .C(_00588_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09932_ (.A1(_03650_),
    .A2(_03653_),
    .B(_03656_),
    .ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09933_ (.A1(_03645_),
    .A2(_03647_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09934_ (.A1(_03568_),
    .A2(_03643_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09935_ (.A1(_03565_),
    .A2(_03644_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09936_ (.A1(_02268_),
    .A2(_02540_),
    .A3(_03639_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09937_ (.A1(_03636_),
    .A2(_03638_),
    .B(_03660_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09938_ (.A1(_03571_),
    .A2(_03632_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09939_ (.A1(_03633_),
    .A2(_03642_),
    .B(_03663_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09940_ (.A1(_03573_),
    .A2(_03604_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09941_ (.A1(_03605_),
    .A2(_03631_),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09942_ (.A1(_03665_),
    .A2(_03666_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09943_ (.A1(_03577_),
    .A2(_03590_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09944_ (.A1(_03591_),
    .A2(_03603_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09945_ (.A1(_03668_),
    .A2(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09946_ (.A1(_02260_),
    .A2(_02386_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09947_ (.A1(_02479_),
    .A2(_02256_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09948_ (.I0(_02387_),
    .I1(_03671_),
    .S(_03673_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09949_ (.A1(_03236_),
    .A2(_02351_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09950_ (.A1(_02263_),
    .A2(_02375_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09951_ (.A1(_02272_),
    .A2(_02655_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09952_ (.A1(_03676_),
    .A2(_03677_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09953_ (.A1(_03675_),
    .A2(_03678_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09954_ (.A1(_03674_),
    .A2(_03679_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09955_ (.A1(_03580_),
    .A2(_03582_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09956_ (.A1(_03583_),
    .A2(_03589_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09957_ (.A1(_03681_),
    .A2(_03682_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09958_ (.A1(_03680_),
    .A2(_03684_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09959_ (.A1(_02277_),
    .A2(_03014_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09960_ (.A1(_03534_),
    .A2(_03686_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09961_ (.A1(_03598_),
    .A2(_03600_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09962_ (.A1(_03687_),
    .A2(_03688_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09963_ (.A1(_03523_),
    .A2(_03676_),
    .B1(_03587_),
    .B2(_03588_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09964_ (.A1(_02296_),
    .A2(_02314_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09965_ (.A1(_02287_),
    .A2(_02326_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09966_ (.A1(_03686_),
    .A2(_03691_),
    .A3(_03692_),
    .Z(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09967_ (.A1(_03690_),
    .A2(_03693_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09968_ (.A1(_03689_),
    .A2(_03695_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09969_ (.A1(_03685_),
    .A2(_03696_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09970_ (.A1(_03670_),
    .A2(_03697_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09971_ (.I(_03698_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09972_ (.A1(_03621_),
    .A2(_03625_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09973_ (.A1(_03617_),
    .A2(_03627_),
    .B(_03700_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09974_ (.A1(_03597_),
    .A2(_03601_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09975_ (.A1(_03594_),
    .A2(_03602_),
    .B(_03702_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09976_ (.A1(_02267_),
    .A2(_02393_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09977_ (.A1(_02433_),
    .A2(_02348_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09978_ (.A1(_02462_),
    .A2(_02359_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09979_ (.A1(_03706_),
    .A2(_03707_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09980_ (.A1(_03704_),
    .A2(_03708_),
    .Z(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09981_ (.A1(_02300_),
    .A2(_03006_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09982_ (.A1(_03504_),
    .A2(_03710_),
    .B1(_03623_),
    .B2(_03624_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09983_ (.A1(_02281_),
    .A2(_02334_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09984_ (.A1(_02290_),
    .A2(_02783_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09985_ (.A1(_03710_),
    .A2(_03713_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09986_ (.A1(_03712_),
    .A2(_03714_),
    .Z(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09987_ (.A1(_03711_),
    .A2(_03715_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09988_ (.A1(_03709_),
    .A2(_03717_),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09989_ (.A1(_03703_),
    .A2(_03718_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09990_ (.A1(_03701_),
    .A2(_03719_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09991_ (.A1(_03699_),
    .A2(_03720_),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09992_ (.A1(_03667_),
    .A2(_03721_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09993_ (.A1(_03612_),
    .A2(_03628_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09994_ (.A1(_03608_),
    .A2(_03630_),
    .B(_03723_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09995_ (.A1(_02282_),
    .A2(_02624_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09996_ (.A1(_03725_),
    .A2(_03706_),
    .B1(_03616_),
    .B2(_03613_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09997_ (.A1(_03724_),
    .A2(_03726_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09998_ (.A1(_02259_),
    .A2(_02539_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09999_ (.A1(_03728_),
    .A2(_03729_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10000_ (.A1(_03722_),
    .A2(_03730_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10001_ (.A1(_03662_),
    .A2(_03664_),
    .A3(_03731_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10002_ (.A1(_03658_),
    .A2(_03659_),
    .B(_03732_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10003_ (.A1(_03658_),
    .A2(_03659_),
    .A3(_03732_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10004_ (.A1(_03733_),
    .A2(_03734_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10005_ (.A1(_03657_),
    .A2(_03652_),
    .B(_03735_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10006_ (.A1(_03657_),
    .A2(_03652_),
    .A3(_03735_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10007_ (.A1(_02152_),
    .A2(_03736_),
    .A3(_03737_),
    .B(_00735_),
    .ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10008_ (.I(_03648_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10009_ (.A1(_03739_),
    .A2(_03735_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10010_ (.A1(_03657_),
    .A2(_03734_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10011_ (.A1(_03649_),
    .A2(_03740_),
    .B(_03741_),
    .C(_03733_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10012_ (.I(_03731_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10013_ (.A1(_03664_),
    .A2(_03743_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10014_ (.A1(_03664_),
    .A2(_03743_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10015_ (.A1(_03662_),
    .A2(_03744_),
    .B(_03745_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10016_ (.A1(_03238_),
    .A2(_02621_),
    .A3(_03678_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10017_ (.A1(_02264_),
    .A2(_02581_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10018_ (.A1(_03586_),
    .A2(_03747_),
    .B(_03749_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10019_ (.A1(_03747_),
    .A2(_03749_),
    .B(_03750_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10020_ (.A1(_03667_),
    .A2(_03721_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10021_ (.A1(_03722_),
    .A2(_03730_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10022_ (.A1(_03752_),
    .A2(_03753_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10023_ (.A1(_03680_),
    .A2(_03684_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10024_ (.A1(_03685_),
    .A2(_03696_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10025_ (.A1(_03755_),
    .A2(_03756_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10026_ (.A1(_02292_),
    .A2(_02310_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10027_ (.A1(_03711_),
    .A2(_03715_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10028_ (.A1(_03709_),
    .A2(_03717_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10029_ (.A1(_03760_),
    .A2(_03761_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10030_ (.A1(_02278_),
    .A2(_02327_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10031_ (.A1(_02435_),
    .A2(_02336_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10032_ (.A1(_02287_),
    .A2(_02315_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10033_ (.A1(_02259_),
    .A2(_02393_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10034_ (.A1(_02961_),
    .A2(_03765_),
    .A3(_03766_),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10035_ (.A1(_03764_),
    .A2(_03767_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10036_ (.A1(_03686_),
    .A2(_03692_),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10037_ (.A1(_03599_),
    .A2(_03763_),
    .B1(_03769_),
    .B2(_03691_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10038_ (.A1(_03763_),
    .A2(_03768_),
    .A3(_03771_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10039_ (.A1(_03758_),
    .A2(_03762_),
    .A3(_03772_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10040_ (.A1(_03757_),
    .A2(_03773_),
    .Z(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10041_ (.A1(_02463_),
    .A2(_02406_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10042_ (.I(_03690_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10043_ (.A1(_03689_),
    .A2(_03695_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10044_ (.A1(_03776_),
    .A2(_03693_),
    .B(_03777_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10045_ (.A1(_02389_),
    .A2(_03673_),
    .B1(_03674_),
    .B2(_03679_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10046_ (.A1(_03775_),
    .A2(_03778_),
    .A3(_03779_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10047_ (.A1(_03622_),
    .A2(_03758_),
    .B1(_03714_),
    .B2(_03712_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10048_ (.A1(_02267_),
    .A2(_02624_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10049_ (.A1(_03238_),
    .A2(_02342_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10050_ (.A1(_03783_),
    .A2(_03784_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10051_ (.A1(_03780_),
    .A2(_03782_),
    .A3(_03785_),
    .Z(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10052_ (.A1(_03703_),
    .A2(_03718_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10053_ (.A1(_03701_),
    .A2(_03719_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10054_ (.A1(_03787_),
    .A2(_03788_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10055_ (.A1(_03615_),
    .A2(_03775_),
    .B1(_03708_),
    .B2(_03704_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10056_ (.A1(_02282_),
    .A2(_02320_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10057_ (.A1(_02273_),
    .A2(_02353_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10058_ (.A1(_02260_),
    .A2(_02377_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10059_ (.A1(_03791_),
    .A2(_03793_),
    .A3(_03794_),
    .Z(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10060_ (.A1(_03789_),
    .A2(_03790_),
    .A3(_03795_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10061_ (.A1(_03774_),
    .A2(_03786_),
    .A3(_03796_),
    .Z(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10062_ (.I(_03724_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10063_ (.A1(_03798_),
    .A2(_03726_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10064_ (.A1(_03728_),
    .A2(_03729_),
    .B(_03799_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10065_ (.A1(_03670_),
    .A2(_03697_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10066_ (.A1(_03699_),
    .A2(_03720_),
    .B(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10067_ (.A1(_03797_),
    .A2(_03800_),
    .A3(_03802_),
    .Z(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10068_ (.A1(_03754_),
    .A2(_03804_),
    .Z(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10069_ (.A1(_03746_),
    .A2(_03751_),
    .A3(_03805_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10070_ (.A1(_03742_),
    .A2(_03806_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10071_ (.A1(_03742_),
    .A2(_03806_),
    .B(_05295_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10072_ (.A1(_03807_),
    .A2(_03808_),
    .B(_00674_),
    .ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10073_ (.I(net31),
    .Z(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10074_ (.I(_03809_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10075_ (.I(_03810_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10076_ (.I(_03811_),
    .Z(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10077_ (.I(_03812_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10078_ (.I(_03814_),
    .Z(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10079_ (.I(_03815_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10080_ (.I(_03816_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10081_ (.I(net30),
    .Z(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10082_ (.I(_03818_),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10083_ (.I(_03819_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10084_ (.I(_03820_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10085_ (.I(net94),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10086_ (.A1(_03821_),
    .A2(_03822_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10087_ (.I(_03821_),
    .Z(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10088_ (.I(net94),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10089_ (.I(_03826_),
    .Z(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10090_ (.A1(_03825_),
    .A2(_03827_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10091_ (.A1(_03817_),
    .A2(_01662_),
    .B1(_01498_),
    .B2(_03823_),
    .C1(_03828_),
    .C2(_01890_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10092_ (.I(_03827_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10093_ (.I(_03830_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10094_ (.I(_03831_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10095_ (.I(_03825_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10096_ (.A1(_03833_),
    .A2(_00734_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10097_ (.I(_03825_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10098_ (.A1(_03836_),
    .A2(_01825_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10099_ (.A1(_03832_),
    .A2(_00950_),
    .B1(_03834_),
    .B2(_03837_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10100_ (.A1(_03829_),
    .A2(_03838_),
    .ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10101_ (.A1(_03833_),
    .A2(_03832_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10102_ (.I(net95),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10103_ (.I(_03840_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10104_ (.I(_03841_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10105_ (.I(_03842_),
    .Z(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10106_ (.A1(_03843_),
    .A2(_03815_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10107_ (.A1(_03839_),
    .A2(_03844_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10108_ (.I(net46),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10109_ (.I(_03847_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10110_ (.I(net110),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10111_ (.A1(_03848_),
    .A2(_03849_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10112_ (.I(net108),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10113_ (.I(_03851_),
    .Z(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10114_ (.I(_03852_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10115_ (.I(net44),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10116_ (.I(_03854_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10117_ (.I(_03855_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10118_ (.A1(_03853_),
    .A2(_03857_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10119_ (.I(net106),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10120_ (.I(_03859_),
    .Z(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10121_ (.I(net42),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10122_ (.I(_03861_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10123_ (.I(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10124_ (.A1(_03860_),
    .A2(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10125_ (.I(net104),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10126_ (.I(_03865_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10127_ (.I(_03866_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10128_ (.I(_03868_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10129_ (.I(_03869_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10130_ (.I(net40),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10131_ (.I(_03871_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10132_ (.I(_03872_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10133_ (.I(_03873_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10134_ (.A1(_03870_),
    .A2(_03874_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10135_ (.A1(_03870_),
    .A2(_03873_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10136_ (.I(net103),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10137_ (.I(_03877_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10138_ (.I(_03879_),
    .Z(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10139_ (.I(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10140_ (.I(net39),
    .Z(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10141_ (.I(_03882_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10142_ (.I(_03883_),
    .Z(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10143_ (.A1(_03881_),
    .A2(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10144_ (.I(net101),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10145_ (.I(_03886_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10146_ (.I(_03887_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10147_ (.I(_03888_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10148_ (.I(_03890_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10149_ (.I(net37),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10150_ (.I(_03892_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10151_ (.I(_03893_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10152_ (.I(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10153_ (.A1(_03891_),
    .A2(_03895_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10154_ (.I(net100),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10155_ (.I(_03897_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10156_ (.I(_03898_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10157_ (.I(_03899_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10158_ (.I(net36),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10159_ (.I(_03902_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10160_ (.I(_03903_),
    .Z(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10161_ (.I(_03904_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10162_ (.A1(_03901_),
    .A2(_03905_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10163_ (.I(net99),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10164_ (.I(_03907_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10165_ (.I(_03908_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10166_ (.I(_03909_),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10167_ (.I(net35),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10168_ (.I(_03912_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10169_ (.I(_03913_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10170_ (.I(_03914_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10171_ (.I(_03915_),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10172_ (.I(_03916_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10173_ (.A1(_03910_),
    .A2(_03917_),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10174_ (.I(net98),
    .Z(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10175_ (.I(net34),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10176_ (.A1(_03919_),
    .A2(_03920_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10177_ (.I(_03919_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10178_ (.I(_03923_),
    .Z(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10179_ (.I(_03924_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10180_ (.I(_03920_),
    .Z(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10181_ (.I(_03926_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10182_ (.I(_03927_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10183_ (.A1(_03925_),
    .A2(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10184_ (.A1(_03921_),
    .A2(_03929_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10185_ (.I(net97),
    .Z(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10186_ (.I(_03931_),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10187_ (.I(_03932_),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10188_ (.I(_03934_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10189_ (.I(_03935_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10190_ (.I(net33),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10191_ (.I(_03937_),
    .Z(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10192_ (.I(_03938_),
    .Z(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10193_ (.I(_03939_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10194_ (.I(_03940_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10195_ (.A1(_03936_),
    .A2(_03941_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10196_ (.I(_03822_),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10197_ (.I(_03814_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10198_ (.I(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10199_ (.A1(_03833_),
    .A2(_03943_),
    .B1(_03843_),
    .B2(_03946_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10200_ (.I(net96),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10201_ (.I(_03948_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10202_ (.I(_03949_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10203_ (.I(_03950_),
    .Z(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10204_ (.I(_03951_),
    .Z(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10205_ (.I(_03952_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10206_ (.I(_03953_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10207_ (.I(net32),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10208_ (.I(_03956_),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10209_ (.I(_03957_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10210_ (.I(_03958_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10211_ (.I(_03959_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10212_ (.I(_03843_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10213_ (.A1(_03954_),
    .A2(_03960_),
    .B1(_03961_),
    .B2(_03946_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10214_ (.A1(_03934_),
    .A2(_03940_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10215_ (.A1(_03931_),
    .A2(_03939_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10216_ (.I(_03964_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10217_ (.A1(_03963_),
    .A2(_03965_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10218_ (.A1(_03954_),
    .A2(_03960_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10219_ (.A1(_03947_),
    .A2(_03962_),
    .B(_03967_),
    .C(_03968_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10220_ (.A1(_03823_),
    .A2(_03844_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10221_ (.A1(_03952_),
    .A2(_03960_),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10222_ (.A1(_03963_),
    .A2(_03965_),
    .B(_03970_),
    .C(_03971_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10223_ (.A1(_03942_),
    .A2(_03969_),
    .B(_03972_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10224_ (.A1(_03909_),
    .A2(_03916_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10225_ (.I(_03925_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10226_ (.I(_03928_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10227_ (.I(_03976_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10228_ (.A1(_03975_),
    .A2(_03978_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10229_ (.A1(_03930_),
    .A2(_03973_),
    .B(_03974_),
    .C(_03979_),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10230_ (.A1(_03901_),
    .A2(_03905_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10231_ (.A1(_03906_),
    .A2(_03918_),
    .A3(_03980_),
    .B(_03981_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10232_ (.A1(_03891_),
    .A2(_03895_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10233_ (.A1(_03881_),
    .A2(_03884_),
    .Z(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10234_ (.A1(_03896_),
    .A2(_03982_),
    .B(_03983_),
    .C(_03984_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10235_ (.A1(_03876_),
    .A2(_03885_),
    .A3(_03985_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10236_ (.I(net105),
    .Z(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10237_ (.I(_03987_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10238_ (.I(_03989_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10239_ (.I(net41),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10240_ (.I(_03991_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10241_ (.A1(_03990_),
    .A2(_03992_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10242_ (.I(_03992_),
    .Z(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10243_ (.A1(_03990_),
    .A2(_03994_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10244_ (.A1(_03993_),
    .A2(_03995_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10245_ (.I(_03996_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10246_ (.I(_03989_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10247_ (.A1(_03998_),
    .A2(_03994_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10248_ (.A1(_03875_),
    .A2(_03986_),
    .A3(_03997_),
    .B(_04000_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10249_ (.A1(_03860_),
    .A2(_03863_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10250_ (.A1(_03864_),
    .A2(_04001_),
    .B(_04002_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10251_ (.I(net107),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10252_ (.I(_04004_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10253_ (.I(_04005_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10254_ (.I(net43),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10255_ (.I(_04007_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10256_ (.I(_04008_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10257_ (.A1(_04006_),
    .A2(_04009_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10258_ (.I(_04006_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10259_ (.A1(_04012_),
    .A2(_04009_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10260_ (.A1(_04003_),
    .A2(_04011_),
    .B(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10261_ (.A1(_03853_),
    .A2(_03857_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10262_ (.A1(_03858_),
    .A2(_04014_),
    .B(_04015_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10263_ (.I(net109),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10264_ (.I(_04017_),
    .Z(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10265_ (.I(net45),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10266_ (.I(_04019_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10267_ (.A1(_04018_),
    .A2(_04020_),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10268_ (.I(_04018_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10269_ (.A1(_04023_),
    .A2(_04020_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10270_ (.A1(_04016_),
    .A2(_04022_),
    .B(_04024_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10271_ (.A1(_03848_),
    .A2(_03849_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10272_ (.A1(_03850_),
    .A2(_04025_),
    .B(_04026_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10273_ (.I(_03894_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10274_ (.A1(_03891_),
    .A2(_04028_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10275_ (.I(_04029_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10276_ (.I(_03930_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10277_ (.A1(_03918_),
    .A2(_03974_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10278_ (.I(_03981_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10279_ (.A1(_03906_),
    .A2(_04034_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10280_ (.A1(_04031_),
    .A2(_04033_),
    .A3(_04035_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10281_ (.A1(_03972_),
    .A2(_04030_),
    .A3(_04036_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10282_ (.I(_04037_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10283_ (.A1(_03852_),
    .A2(_03855_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10284_ (.I(_03860_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10285_ (.I(_03862_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10286_ (.A1(_04040_),
    .A2(_04041_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10287_ (.A1(_03869_),
    .A2(_03874_),
    .Z(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10288_ (.A1(_04022_),
    .A2(_04039_),
    .A3(_04042_),
    .A4(_04044_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10289_ (.I(_03984_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10290_ (.I(_03996_),
    .Z(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10291_ (.I(_04009_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10292_ (.A1(_04012_),
    .A2(_04048_),
    .Z(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10293_ (.A1(_03850_),
    .A2(_04046_),
    .A3(_04047_),
    .A4(_04049_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10294_ (.A1(_04038_),
    .A2(_04045_),
    .A3(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10295_ (.A1(_04027_),
    .A2(_04051_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10296_ (.I(_04052_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10297_ (.I(_04053_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10298_ (.A1(_03823_),
    .A2(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10299_ (.A1(_03846_),
    .A2(_04056_),
    .B(_04756_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10300_ (.A1(_03846_),
    .A2(_04056_),
    .B(_04057_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10301_ (.A1(_03836_),
    .A2(_03830_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10302_ (.I(_03961_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10303_ (.I(_04060_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10304_ (.A1(_04061_),
    .A2(_03817_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10305_ (.A1(_04059_),
    .A2(_04062_),
    .B(_00045_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10306_ (.A1(_04059_),
    .A2(_04062_),
    .B(_04063_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10307_ (.I(_03959_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _10308_ (.A1(_04066_),
    .A2(_00233_),
    .B1(_00414_),
    .B2(_03946_),
    .C1(_04269_),
    .C2(_03836_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10309_ (.A1(_04571_),
    .A2(_04061_),
    .B(_04062_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10310_ (.A1(_03836_),
    .A2(_04060_),
    .B1(_03817_),
    .B2(_03832_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10311_ (.A1(_03961_),
    .A2(_03816_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10312_ (.A1(_04059_),
    .A2(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10313_ (.A1(_00951_),
    .A2(_04069_),
    .A3(_04071_),
    .B1(_00959_),
    .B2(_04070_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10314_ (.A1(_04060_),
    .A2(_00421_),
    .B1(_04068_),
    .B2(_04604_),
    .C(_04072_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10315_ (.A1(_04058_),
    .A2(_04064_),
    .A3(_04067_),
    .A4(_04073_),
    .ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10316_ (.I(_03971_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10317_ (.A1(_03961_),
    .A2(_03816_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10318_ (.A1(_03828_),
    .A2(_03844_),
    .B(_04076_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10319_ (.A1(_04074_),
    .A2(_04077_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10320_ (.A1(_02495_),
    .A2(_04078_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10321_ (.I(_03941_),
    .Z(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10322_ (.A1(_03953_),
    .A2(_03959_),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10323_ (.A1(_04080_),
    .A2(_00211_),
    .B1(_04204_),
    .B2(_04081_),
    .C1(_00212_),
    .C2(_03817_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10324_ (.A1(_04066_),
    .A2(_00734_),
    .B1(_04074_),
    .B2(_04388_),
    .C(_04082_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10325_ (.A1(_03954_),
    .A2(_00950_),
    .B(_04083_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10326_ (.A1(_03823_),
    .A2(_03844_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10327_ (.I(_04053_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10328_ (.A1(_03839_),
    .A2(_04062_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10329_ (.A1(_04060_),
    .A2(_03946_),
    .B(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10330_ (.A1(_04074_),
    .A2(_04089_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10331_ (.A1(_04085_),
    .A2(_04087_),
    .A3(_04090_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10332_ (.A1(_04085_),
    .A2(_04087_),
    .B(_04090_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10333_ (.A1(_03254_),
    .A2(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10334_ (.A1(_03820_),
    .A2(_03951_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10335_ (.A1(_04076_),
    .A2(_04094_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10336_ (.I(_03827_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10337_ (.A1(_04096_),
    .A2(_04066_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10338_ (.A1(_04095_),
    .A2(_04098_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10339_ (.A1(_04095_),
    .A2(_04098_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10340_ (.A1(_04071_),
    .A2(_04099_),
    .A3(_04100_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10341_ (.A1(_04099_),
    .A2(_04100_),
    .B(_04071_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10342_ (.A1(_00992_),
    .A2(_04102_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10343_ (.A1(_04091_),
    .A2(_04093_),
    .B1(_04101_),
    .B2(_04103_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10344_ (.A1(_04079_),
    .A2(_04084_),
    .A3(_04104_),
    .ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10345_ (.A1(_03947_),
    .A2(_03962_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10346_ (.A1(_03954_),
    .A2(_03960_),
    .B(_04105_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10347_ (.I(_04052_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10348_ (.A1(_04074_),
    .A2(_04089_),
    .B(_04053_),
    .C(_03968_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10349_ (.A1(_04106_),
    .A2(_04108_),
    .B(_04109_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10350_ (.A1(_03967_),
    .A2(_04110_),
    .Z(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10351_ (.A1(_03952_),
    .A2(_03815_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10352_ (.A1(_03959_),
    .A2(_03842_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10353_ (.A1(_03825_),
    .A2(_03935_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10354_ (.A1(_04112_),
    .A2(_04113_),
    .A3(_04114_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10355_ (.A1(_03821_),
    .A2(_03953_),
    .A3(_03843_),
    .A4(_03815_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10356_ (.A1(_03826_),
    .A2(_03941_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10357_ (.A1(_04116_),
    .A2(_04117_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10358_ (.A1(_04115_),
    .A2(_04119_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10359_ (.A1(_04099_),
    .A2(_04101_),
    .Z(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10360_ (.A1(_04120_),
    .A2(_04121_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10361_ (.I(_03949_),
    .Z(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10362_ (.A1(_04123_),
    .A2(_03958_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10363_ (.A1(_03971_),
    .A2(_04077_),
    .B(_04124_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10364_ (.A1(_03967_),
    .A2(_04125_),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10365_ (.I(_03965_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10366_ (.A1(_00395_),
    .A2(_04127_),
    .B(_03963_),
    .C(_04366_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10367_ (.A1(_03976_),
    .A2(_05191_),
    .B1(_05267_),
    .B2(_04066_),
    .C(_04128_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10368_ (.A1(_03935_),
    .A2(_00240_),
    .B1(_04127_),
    .B2(_01035_),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10369_ (.A1(_04080_),
    .A2(_01238_),
    .B(_04130_),
    .C(_04131_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10370_ (.A1(_00244_),
    .A2(_04122_),
    .B1(_04126_),
    .B2(_02580_),
    .C(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10371_ (.A1(_00762_),
    .A2(_04111_),
    .B(_04133_),
    .ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10372_ (.I(_04027_),
    .Z(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10373_ (.A1(_04031_),
    .A2(_03973_),
    .Z(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10374_ (.A1(_03972_),
    .A2(_04134_),
    .B(_04135_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10375_ (.A1(_03972_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10376_ (.A1(_05292_),
    .A2(_04137_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10377_ (.A1(_03935_),
    .A2(_04080_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10378_ (.A1(_04140_),
    .A2(_04125_),
    .B(_04127_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10379_ (.A1(_04031_),
    .A2(_04141_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10380_ (.I(_03921_),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10381_ (.A1(_05202_),
    .A2(_04143_),
    .B(_03929_),
    .C(_00397_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10382_ (.A1(_03915_),
    .A2(_00130_),
    .B1(_00394_),
    .B2(_04080_),
    .C(_04144_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10383_ (.A1(_03975_),
    .A2(_05583_),
    .B1(_04143_),
    .B2(_02692_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10384_ (.A1(_03976_),
    .A2(_05180_),
    .B(_04145_),
    .C(_04146_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10385_ (.A1(_04485_),
    .A2(_04142_),
    .B(_04147_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10386_ (.A1(_04099_),
    .A2(_04120_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10387_ (.A1(_04101_),
    .A2(_04120_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10388_ (.A1(_04116_),
    .A2(_04117_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10389_ (.A1(_04115_),
    .A2(_04119_),
    .B(_04152_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10390_ (.A1(_03819_),
    .A2(_03924_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10391_ (.A1(_03932_),
    .A2(_03812_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10392_ (.A1(_03940_),
    .A2(_03842_),
    .Z(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10393_ (.A1(_04124_),
    .A2(_04155_),
    .A3(_04156_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10394_ (.A1(_04154_),
    .A2(_04157_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10395_ (.A1(_03820_),
    .A2(_03932_),
    .B1(_03951_),
    .B2(_03814_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10396_ (.A1(_04094_),
    .A2(_04155_),
    .B1(_04159_),
    .B2(_04113_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10397_ (.A1(_03822_),
    .A2(_03927_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10398_ (.A1(_04160_),
    .A2(_04162_),
    .Z(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10399_ (.A1(_04153_),
    .A2(_04158_),
    .A3(_04163_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10400_ (.A1(_04149_),
    .A2(_04151_),
    .A3(_04164_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10401_ (.A1(_02152_),
    .A2(_04165_),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10402_ (.A1(_04136_),
    .A2(_04138_),
    .B(_04148_),
    .C(_04166_),
    .ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10403_ (.A1(_04031_),
    .A2(_03973_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10404_ (.I(_04052_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10405_ (.A1(_03975_),
    .A2(_03978_),
    .B(_03942_),
    .C(_03969_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10406_ (.A1(_03979_),
    .A2(_04169_),
    .B(_04053_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10407_ (.A1(_03979_),
    .A2(_04167_),
    .A3(_04168_),
    .B(_04170_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10408_ (.A1(_04033_),
    .A2(_04172_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10409_ (.A1(_04149_),
    .A2(_04164_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10410_ (.A1(_04149_),
    .A2(_04164_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10411_ (.A1(_04151_),
    .A2(_04174_),
    .B(_04175_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10412_ (.A1(_04158_),
    .A2(_04163_),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10413_ (.A1(_04153_),
    .A2(_04177_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10414_ (.A1(_03943_),
    .A2(_03928_),
    .A3(_04160_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10415_ (.A1(_04158_),
    .A2(_04163_),
    .B(_04179_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10416_ (.A1(_04124_),
    .A2(_04155_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10417_ (.I(_03931_),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10418_ (.A1(_04183_),
    .A2(_03957_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10419_ (.A1(_04112_),
    .A2(_04184_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10420_ (.A1(_04156_),
    .A2(_04181_),
    .B(_04185_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10421_ (.A1(_03822_),
    .A2(_03915_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10422_ (.A1(_04186_),
    .A2(_04187_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10423_ (.A1(_03821_),
    .A2(_03925_),
    .A3(_04157_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10424_ (.I(net30),
    .Z(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10425_ (.I(_04190_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10426_ (.I(net99),
    .Z(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10427_ (.I(_04192_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10428_ (.I(_04194_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10429_ (.A1(_04191_),
    .A2(_04195_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10430_ (.A1(_03925_),
    .A2(_03814_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10431_ (.A1(_03820_),
    .A2(_03909_),
    .A3(_03924_),
    .A4(_03812_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10432_ (.A1(_04196_),
    .A2(_04197_),
    .B(_04198_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10433_ (.A1(_03926_),
    .A2(_03841_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10434_ (.A1(_03940_),
    .A2(_03951_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10435_ (.A1(_04184_),
    .A2(_04200_),
    .A3(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10436_ (.A1(_04199_),
    .A2(_04202_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10437_ (.A1(_04189_),
    .A2(_04203_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10438_ (.A1(_04180_),
    .A2(_04188_),
    .A3(_04205_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10439_ (.A1(_04178_),
    .A2(_04206_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10440_ (.A1(_04176_),
    .A2(_04207_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10441_ (.A1(_03930_),
    .A2(_04141_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10442_ (.I(_04033_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10443_ (.A1(_04143_),
    .A2(_04209_),
    .B(_04210_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10444_ (.A1(_04143_),
    .A2(_04210_),
    .A3(_04209_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10445_ (.A1(_01423_),
    .A2(_04212_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10446_ (.I(net35),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10447_ (.A1(_04192_),
    .A2(_04214_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10448_ (.I(_04216_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10449_ (.I(_03905_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _10450_ (.A1(_04218_),
    .A2(_00232_),
    .B1(_00131_),
    .B2(_03917_),
    .C1(_04258_),
    .C2(_03976_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10451_ (.A1(_04388_),
    .A2(_04033_),
    .B1(_04217_),
    .B2(_00959_),
    .C(_04219_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10452_ (.A1(_03910_),
    .A2(_02744_),
    .B1(_04211_),
    .B2(_04213_),
    .C(_04220_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10453_ (.A1(_00137_),
    .A2(_04173_),
    .B1(_04208_),
    .B2(_02812_),
    .C(_04221_),
    .ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10454_ (.A1(_04188_),
    .A2(_04205_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10455_ (.A1(_04180_),
    .A2(_04222_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10456_ (.A1(_04178_),
    .A2(_04206_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10457_ (.A1(_04176_),
    .A2(_04207_),
    .B(_04224_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10458_ (.A1(_04199_),
    .A2(_04202_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10459_ (.A1(_03913_),
    .A2(_03841_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10460_ (.A1(_03927_),
    .A2(_04123_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10461_ (.A1(_03964_),
    .A2(_04228_),
    .A3(_04229_),
    .Z(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10462_ (.I(_03809_),
    .Z(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10463_ (.A1(_03908_),
    .A2(_04231_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10464_ (.A1(_03923_),
    .A2(_03957_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10465_ (.I(net100),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10466_ (.I(_04234_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10467_ (.I(_04235_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10468_ (.A1(_03819_),
    .A2(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10469_ (.A1(_04232_),
    .A2(_04233_),
    .A3(_04238_),
    .Z(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10470_ (.A1(_04198_),
    .A2(_04230_),
    .A3(_04239_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10471_ (.A1(_04227_),
    .A2(_04240_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10472_ (.A1(_04189_),
    .A2(_04203_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10473_ (.A1(_03943_),
    .A2(_03905_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10474_ (.I(_04200_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10475_ (.A1(_04184_),
    .A2(_04201_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10476_ (.A1(_04081_),
    .A2(_04127_),
    .B1(_04244_),
    .B2(_04245_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10477_ (.A1(_04242_),
    .A2(_04243_),
    .A3(_04246_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10478_ (.A1(_04186_),
    .A2(_04187_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10479_ (.A1(_04188_),
    .A2(_04205_),
    .B(_04249_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10480_ (.A1(_04241_),
    .A2(_04248_),
    .A3(_04250_),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10481_ (.A1(_04223_),
    .A2(_04226_),
    .A3(_04251_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10482_ (.I(_04035_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10483_ (.A1(_04253_),
    .A2(_04211_),
    .A3(_04217_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10484_ (.A1(_04211_),
    .A2(_04217_),
    .B(_04035_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10485_ (.A1(_04254_),
    .A2(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10486_ (.I(net36),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10487_ (.A1(_03897_),
    .A2(_04257_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10488_ (.A1(_03917_),
    .A2(_01858_),
    .A3(_04065_),
    .B1(_04615_),
    .B2(_04218_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10489_ (.A1(_04028_),
    .A2(_00232_),
    .B1(_04204_),
    .B2(_04259_),
    .C(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10490_ (.A1(_04218_),
    .A2(_02822_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10491_ (.A1(_01379_),
    .A2(_04253_),
    .B(_04261_),
    .C(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10492_ (.A1(_03899_),
    .A2(_05498_),
    .B1(_04256_),
    .B2(_05503_),
    .C(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10493_ (.I(_04027_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10494_ (.A1(_03910_),
    .A2(_03917_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10495_ (.A1(_03974_),
    .A2(_03979_),
    .A3(_04169_),
    .B(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10496_ (.A1(_04265_),
    .A2(_04051_),
    .B(_04267_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10497_ (.A1(_03918_),
    .A2(_03980_),
    .A3(_04108_),
    .B(_04268_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10498_ (.I(_01477_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10499_ (.A1(_04253_),
    .A2(_04270_),
    .B(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10500_ (.A1(_04253_),
    .A2(_04270_),
    .B(_04272_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10501_ (.A1(_02977_),
    .A2(_04252_),
    .B(_04264_),
    .C(_04273_),
    .ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10502_ (.A1(_03981_),
    .A2(_04267_),
    .B(_03906_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10503_ (.A1(_03982_),
    .A2(_04168_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10504_ (.A1(_04168_),
    .A2(_04274_),
    .B(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10505_ (.A1(_04030_),
    .A2(_04276_),
    .Z(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10506_ (.I(_04241_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10507_ (.A1(_04278_),
    .A2(_04248_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10508_ (.A1(_04280_),
    .A2(_04250_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10509_ (.A1(_04223_),
    .A2(_04251_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10510_ (.A1(_04223_),
    .A2(_04251_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10511_ (.A1(_04226_),
    .A2(_04282_),
    .B(_04283_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10512_ (.A1(_04278_),
    .A2(_04248_),
    .Z(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10513_ (.A1(_04242_),
    .A2(_04246_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10514_ (.A1(_04242_),
    .A2(_04246_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10515_ (.A1(_04243_),
    .A2(_04286_),
    .B(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10516_ (.A1(_03819_),
    .A2(_03888_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10517_ (.A1(_04154_),
    .A2(_04232_),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10518_ (.A1(_04291_),
    .A2(_04239_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10519_ (.A1(_04291_),
    .A2(_04239_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10520_ (.A1(_04230_),
    .A2(_04292_),
    .B(_04293_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10521_ (.I(_03840_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10522_ (.A1(_03904_),
    .A2(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10523_ (.I(net97),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10524_ (.A1(_03920_),
    .A2(_04297_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10525_ (.A1(_03913_),
    .A2(_03949_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10526_ (.A1(_04298_),
    .A2(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10527_ (.A1(_04296_),
    .A2(_04300_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10528_ (.A1(_03897_),
    .A2(_03809_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10529_ (.A1(_03818_),
    .A2(_04237_),
    .B1(_04195_),
    .B2(_03811_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10530_ (.A1(_04196_),
    .A2(_04303_),
    .B1(_04304_),
    .B2(_04233_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10531_ (.I(net98),
    .Z(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10532_ (.I(net33),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10533_ (.A1(_04306_),
    .A2(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10534_ (.I(_03956_),
    .Z(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10535_ (.A1(_04194_),
    .A2(_04309_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10536_ (.A1(_04303_),
    .A2(_04308_),
    .A3(_04310_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10537_ (.A1(_04305_),
    .A2(_04311_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10538_ (.A1(_04302_),
    .A2(_04313_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10539_ (.I(_04314_),
    .Z(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10540_ (.A1(_04289_),
    .A2(_04294_),
    .A3(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10541_ (.A1(_03827_),
    .A2(_03894_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10542_ (.A1(_04227_),
    .A2(_04240_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10543_ (.A1(_03927_),
    .A2(_03953_),
    .B(_03965_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10544_ (.A1(_04228_),
    .A2(_04319_),
    .B1(_04298_),
    .B2(_04201_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10545_ (.A1(_04318_),
    .A2(_04320_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10546_ (.A1(_04316_),
    .A2(_04317_),
    .A3(_04321_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10547_ (.A1(_04285_),
    .A2(_04288_),
    .A3(_04322_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10548_ (.A1(_04281_),
    .A2(_04284_),
    .A3(_04324_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10549_ (.A1(_04030_),
    .A2(_04255_),
    .A3(_04259_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10550_ (.A1(_04255_),
    .A2(_04259_),
    .B(_04029_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10551_ (.A1(_04326_),
    .A2(_04327_),
    .Z(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10552_ (.I(net37),
    .Z(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10553_ (.A1(_03886_),
    .A2(_04329_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10554_ (.I(_04330_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10555_ (.I(_04331_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10556_ (.A1(_04218_),
    .A2(_01073_),
    .B1(_04332_),
    .B2(_01577_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10557_ (.I(_03884_),
    .Z(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10558_ (.A1(_04335_),
    .A2(_01417_),
    .B1(_05505_),
    .B2(_03895_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10559_ (.A1(_04028_),
    .A2(_05586_),
    .B1(_00133_),
    .B2(_04030_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10560_ (.A1(_04333_),
    .A2(_04336_),
    .A3(_04337_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10561_ (.A1(_03891_),
    .A2(_02744_),
    .B1(_04328_),
    .B2(_02751_),
    .C(_04338_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10562_ (.A1(_00137_),
    .A2(_04277_),
    .B1(_04325_),
    .B2(_02812_),
    .C(_04339_),
    .ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10563_ (.A1(_04281_),
    .A2(_04324_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10564_ (.A1(_04281_),
    .A2(_04324_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10565_ (.A1(_04284_),
    .A2(_04340_),
    .B(_04341_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10566_ (.A1(_04285_),
    .A2(_04322_),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10567_ (.A1(_04285_),
    .A2(_04322_),
    .Z(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10568_ (.A1(_04288_),
    .A2(_04343_),
    .B(_04345_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10569_ (.A1(_04317_),
    .A2(_04321_),
    .Z(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10570_ (.A1(_04316_),
    .A2(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10571_ (.A1(_04317_),
    .A2(_04321_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10572_ (.A1(_04318_),
    .A2(_04320_),
    .B(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10573_ (.I(_04294_),
    .Z(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10574_ (.A1(_04351_),
    .A2(_04314_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10575_ (.A1(_04351_),
    .A2(_04315_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10576_ (.A1(_04289_),
    .A2(_04352_),
    .A3(_04353_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10577_ (.A1(_03826_),
    .A2(_03883_),
    .Z(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10578_ (.A1(_04298_),
    .A2(_04299_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10579_ (.A1(_04296_),
    .A2(_04300_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10580_ (.A1(_04357_),
    .A2(_04358_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10581_ (.A1(_04352_),
    .A2(_04356_),
    .A3(_04359_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10582_ (.A1(_04191_),
    .A2(_03879_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10583_ (.A1(_03890_),
    .A2(_03816_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10584_ (.A1(_03877_),
    .A2(_04231_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10585_ (.A1(_04289_),
    .A2(_04363_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10586_ (.A1(_04361_),
    .A2(_04362_),
    .B(_04364_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10587_ (.A1(_04305_),
    .A2(_04311_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10588_ (.A1(_04302_),
    .A2(_04313_),
    .B(_04367_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10589_ (.A1(_03893_),
    .A2(_04295_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10590_ (.A1(_03903_),
    .A2(_03914_),
    .A3(_04183_),
    .A4(_03950_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10591_ (.A1(_03914_),
    .A2(_04183_),
    .B1(_04123_),
    .B2(_03903_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10592_ (.A1(_04370_),
    .A2(_04371_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10593_ (.A1(_04369_),
    .A2(_04372_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10594_ (.I(_03897_),
    .Z(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10595_ (.I(_03956_),
    .Z(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10596_ (.A1(_04374_),
    .A2(_04375_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10597_ (.A1(_03909_),
    .A2(_03958_),
    .B1(_03812_),
    .B2(_03899_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10598_ (.A1(_04232_),
    .A2(_04376_),
    .B1(_04378_),
    .B2(_04308_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10599_ (.A1(_04195_),
    .A2(_03939_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10600_ (.A1(_03921_),
    .A2(_04376_),
    .A3(_04380_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10601_ (.A1(_04379_),
    .A2(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10602_ (.A1(_04373_),
    .A2(_04382_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10603_ (.A1(_04368_),
    .A2(_04383_),
    .Z(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10604_ (.A1(_04365_),
    .A2(_04384_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10605_ (.A1(_04354_),
    .A2(_04360_),
    .A3(_04385_),
    .Z(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10606_ (.A1(_04348_),
    .A2(_04350_),
    .A3(_04386_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10607_ (.A1(_04342_),
    .A2(_04346_),
    .A3(_04387_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10608_ (.A1(_04046_),
    .A2(_04327_),
    .A3(_04331_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10609_ (.A1(_04327_),
    .A2(_04331_),
    .B(_04046_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10610_ (.A1(_00964_),
    .A2(_04391_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10611_ (.I(net39),
    .Z(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10612_ (.A1(net103),
    .A2(_04393_),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10613_ (.I(_04394_),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10614_ (.A1(_00418_),
    .A2(_04395_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10615_ (.A1(_03880_),
    .A2(_04335_),
    .B(_01123_),
    .C(_04396_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10616_ (.A1(_03880_),
    .A2(_00988_),
    .B1(_04395_),
    .B2(_00989_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10617_ (.I(_03874_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10618_ (.A1(_04335_),
    .A2(_04279_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10619_ (.A1(_04400_),
    .A2(_01651_),
    .B1(_00126_),
    .B2(_04028_),
    .C(_04401_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10620_ (.A1(_04397_),
    .A2(_04398_),
    .A3(_04402_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10621_ (.A1(_04390_),
    .A2(_04392_),
    .B(_04403_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10622_ (.A1(_03896_),
    .A2(_03982_),
    .B(_03983_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10623_ (.A1(_04046_),
    .A2(_04405_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10624_ (.A1(_04134_),
    .A2(_04038_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10625_ (.A1(_04406_),
    .A2(_04407_),
    .B(_04271_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10626_ (.A1(_04406_),
    .A2(_04407_),
    .B(_04408_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10627_ (.A1(_00675_),
    .A2(_04389_),
    .B(_04404_),
    .C(_04409_),
    .ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10628_ (.A1(_04346_),
    .A2(_04387_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10629_ (.A1(_04346_),
    .A2(_04387_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10630_ (.A1(_04342_),
    .A2(_04411_),
    .B(_04412_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10631_ (.A1(_04316_),
    .A2(_04347_),
    .A3(_04386_),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10632_ (.A1(_04316_),
    .A2(_04347_),
    .B(_04386_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10633_ (.A1(_04350_),
    .A2(_04414_),
    .A3(_04415_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10634_ (.A1(_04351_),
    .A2(_04315_),
    .B(_04359_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10635_ (.A1(_04351_),
    .A2(_04315_),
    .A3(_04359_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10636_ (.A1(_04356_),
    .A2(_04417_),
    .B(_04418_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10637_ (.I(_04419_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10638_ (.A1(_04354_),
    .A2(_04385_),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10639_ (.A1(_04354_),
    .A2(_04385_),
    .Z(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10640_ (.A1(_04360_),
    .A2(_04422_),
    .B(_04423_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10641_ (.A1(_04365_),
    .A2(_04384_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10642_ (.A1(_03887_),
    .A2(_03957_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10643_ (.A1(_04191_),
    .A2(_03868_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10644_ (.A1(_04363_),
    .A2(_04426_),
    .A3(_04427_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10645_ (.A1(_04364_),
    .A2(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10646_ (.A1(_04379_),
    .A2(_04381_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10647_ (.A1(_04373_),
    .A2(_04382_),
    .B(_04430_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10648_ (.I(_04257_),
    .Z(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10649_ (.A1(_04433_),
    .A2(_03931_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10650_ (.A1(_03882_),
    .A2(_03840_),
    .Z(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10651_ (.A1(_03893_),
    .A2(_03950_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10652_ (.A1(_04434_),
    .A2(_04435_),
    .A3(_04436_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10653_ (.A1(_04234_),
    .A2(_03937_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10654_ (.I(_04192_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10655_ (.A1(_04439_),
    .A2(_03938_),
    .B1(_04375_),
    .B2(_03898_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10656_ (.I(net34),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10657_ (.A1(_03919_),
    .A2(_04441_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10658_ (.A1(_04310_),
    .A2(_04438_),
    .B1(_04440_),
    .B2(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10659_ (.A1(_03912_),
    .A2(net98),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10660_ (.I(net34),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10661_ (.A1(_04192_),
    .A2(_04446_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10662_ (.A1(_04438_),
    .A2(_04445_),
    .A3(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10663_ (.A1(_04444_),
    .A2(_04448_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10664_ (.A1(_04437_),
    .A2(_04449_),
    .Z(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10665_ (.A1(_04429_),
    .A2(_04432_),
    .A3(_04450_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10666_ (.A1(_04368_),
    .A2(_04383_),
    .Z(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10667_ (.A1(_03943_),
    .A2(_03873_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10668_ (.A1(_04369_),
    .A2(_04372_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10669_ (.A1(_04370_),
    .A2(_04455_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10670_ (.A1(_04452_),
    .A2(_04454_),
    .A3(_04456_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10671_ (.A1(_04425_),
    .A2(_04451_),
    .A3(_04457_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10672_ (.A1(_04421_),
    .A2(_04424_),
    .A3(_04458_),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10673_ (.A1(_04414_),
    .A2(_04416_),
    .B(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10674_ (.I(_04460_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10675_ (.A1(_04414_),
    .A2(_04416_),
    .A3(_04459_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10676_ (.A1(_04461_),
    .A2(_04462_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10677_ (.A1(_04413_),
    .A2(_04463_),
    .Z(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10678_ (.I(_04044_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10679_ (.A1(_04395_),
    .A2(_04466_),
    .A3(_04391_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10680_ (.A1(_04395_),
    .A2(_04391_),
    .B(_04044_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10681_ (.A1(_04467_),
    .A2(_04468_),
    .Z(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10682_ (.I(_03994_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10683_ (.A1(_03869_),
    .A2(_03873_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10684_ (.I(_04471_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10685_ (.A1(_04400_),
    .A2(_00049_),
    .B1(_05591_),
    .B2(_04472_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10686_ (.A1(_04470_),
    .A2(_05511_),
    .B1(_01073_),
    .B2(_04335_),
    .C(_04473_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10687_ (.A1(_04400_),
    .A2(_01265_),
    .B1(_05585_),
    .B2(_04466_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10688_ (.A1(_04474_),
    .A2(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10689_ (.A1(_03869_),
    .A2(_05498_),
    .B1(_04469_),
    .B2(_05503_),
    .C(_04476_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10690_ (.A1(_03885_),
    .A2(_03985_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10691_ (.I(_04051_),
    .Z(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10692_ (.A1(_03881_),
    .A2(_03884_),
    .B1(_03896_),
    .B2(_04274_),
    .C(_03983_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10693_ (.A1(_03885_),
    .A2(_04480_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10694_ (.A1(_04265_),
    .A2(_04479_),
    .B(_04481_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10695_ (.A1(_04478_),
    .A2(_04087_),
    .B(_04482_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10696_ (.A1(_04466_),
    .A2(_04483_),
    .B(_04271_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10697_ (.A1(_04466_),
    .A2(_04483_),
    .B(_04484_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10698_ (.A1(_00675_),
    .A2(_04465_),
    .B(_04477_),
    .C(_04486_),
    .ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10699_ (.I(_04047_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10700_ (.A1(_03876_),
    .A2(_03885_),
    .A3(_04480_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10701_ (.A1(_03870_),
    .A2(_03874_),
    .B(_04488_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10702_ (.A1(_04134_),
    .A2(_04479_),
    .B(_04489_),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10703_ (.A1(_03875_),
    .A2(_03986_),
    .A3(_04055_),
    .B(_04490_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10704_ (.A1(_04487_),
    .A2(_04491_),
    .B(_03254_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10705_ (.A1(_04487_),
    .A2(_04491_),
    .B(_04492_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10706_ (.A1(_04424_),
    .A2(_04458_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10707_ (.A1(_04424_),
    .A2(_04458_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10708_ (.A1(_04421_),
    .A2(_04494_),
    .B(_04496_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10709_ (.A1(_04370_),
    .A2(_04455_),
    .A3(_04452_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10710_ (.A1(_04370_),
    .A2(_04455_),
    .B(_04452_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10711_ (.A1(_04454_),
    .A2(_04498_),
    .B(_04499_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10712_ (.A1(_04365_),
    .A2(_04384_),
    .B(_04451_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10713_ (.A1(_04365_),
    .A2(_04384_),
    .A3(_04451_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10714_ (.A1(_04501_),
    .A2(_04457_),
    .B(_04502_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10715_ (.A1(_04432_),
    .A2(_04450_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10716_ (.A1(_04429_),
    .A2(_04504_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10717_ (.A1(_03818_),
    .A2(_03987_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10718_ (.A1(_03865_),
    .A2(_03810_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10719_ (.A1(_03818_),
    .A2(_03866_),
    .B1(_03877_),
    .B2(_03811_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10720_ (.A1(_04361_),
    .A2(_04508_),
    .B1(_04509_),
    .B2(_04426_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10721_ (.A1(_03886_),
    .A2(_04307_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10722_ (.I(net103),
    .Z(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10723_ (.A1(_04512_),
    .A2(_04309_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10724_ (.A1(_04508_),
    .A2(_04511_),
    .A3(_04513_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10725_ (.A1(_04510_),
    .A2(_04514_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10726_ (.A1(_04507_),
    .A2(_04515_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10727_ (.I(_04516_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10728_ (.A1(_04364_),
    .A2(_04428_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10729_ (.A1(_04444_),
    .A2(_04448_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10730_ (.A1(_04437_),
    .A2(_04449_),
    .B(_04520_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10731_ (.A1(_03892_),
    .A2(_04297_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10732_ (.A1(_03871_),
    .A2(_03840_),
    .Z(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10733_ (.A1(_03882_),
    .A2(_03949_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10734_ (.A1(_04522_),
    .A2(_04523_),
    .A3(_04524_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10735_ (.A1(_04374_),
    .A2(_04441_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10736_ (.A1(_03908_),
    .A2(_03926_),
    .B1(_03939_),
    .B2(_04237_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10737_ (.A1(_04380_),
    .A2(_04526_),
    .B1(_04527_),
    .B2(_04445_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10738_ (.A1(_03902_),
    .A2(_03919_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10739_ (.A1(_04217_),
    .A2(_04526_),
    .A3(_04530_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10740_ (.A1(_04525_),
    .A2(_04529_),
    .A3(_04531_),
    .Z(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10741_ (.A1(_04519_),
    .A2(_04521_),
    .A3(_04532_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10742_ (.A1(_04518_),
    .A2(_04533_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10743_ (.A1(_04432_),
    .A2(_04450_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10744_ (.A1(_03826_),
    .A2(_03991_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10745_ (.A1(_04434_),
    .A2(_04436_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10746_ (.A1(_04434_),
    .A2(_04436_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10747_ (.A1(_04435_),
    .A2(_04537_),
    .B(_04538_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10748_ (.A1(_04535_),
    .A2(_04536_),
    .A3(_04540_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10749_ (.A1(_04505_),
    .A2(_04534_),
    .A3(_04541_),
    .Z(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10750_ (.A1(_04503_),
    .A2(_04542_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10751_ (.A1(_04500_),
    .A2(_04543_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10752_ (.A1(_04497_),
    .A2(_04544_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10753_ (.A1(_04413_),
    .A2(_04462_),
    .B(_04460_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10754_ (.A1(_04545_),
    .A2(_04546_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10755_ (.A1(_04487_),
    .A2(_04468_),
    .A3(_04472_),
    .Z(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10756_ (.A1(_04468_),
    .A2(_04472_),
    .B(_04047_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10757_ (.A1(_04548_),
    .A2(_04549_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10758_ (.I(_04041_),
    .Z(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10759_ (.A1(_04470_),
    .A2(_04279_),
    .B1(_05321_),
    .B2(_04487_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10760_ (.A1(_04552_),
    .A2(_01338_),
    .B1(_03993_),
    .B2(_05320_),
    .C(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10761_ (.A1(_03990_),
    .A2(_04470_),
    .Z(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10762_ (.A1(_03990_),
    .A2(_01493_),
    .B1(_00984_),
    .B2(_04400_),
    .C1(_04555_),
    .C2(_01263_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10763_ (.A1(_04554_),
    .A2(_04556_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10764_ (.A1(_01430_),
    .A2(_04547_),
    .B1(_04551_),
    .B2(_02495_),
    .C(_04557_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10765_ (.A1(_04493_),
    .A2(_04558_),
    .ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10766_ (.I(_04042_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10767_ (.A1(_03998_),
    .A2(_03994_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10768_ (.A1(_04047_),
    .A2(_04489_),
    .B(_04561_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10769_ (.A1(_04001_),
    .A2(_04168_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10770_ (.A1(_04108_),
    .A2(_04562_),
    .B(_04563_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10771_ (.A1(_04559_),
    .A2(_04564_),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10772_ (.I(_04497_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10773_ (.A1(_04566_),
    .A2(_04544_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10774_ (.A1(_04545_),
    .A2(_04546_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10775_ (.A1(_04567_),
    .A2(_04568_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10776_ (.A1(_04503_),
    .A2(_04542_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10777_ (.A1(_04500_),
    .A2(_04543_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10778_ (.A1(_04570_),
    .A2(_04572_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10779_ (.A1(_04535_),
    .A2(_04540_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10780_ (.A1(_04535_),
    .A2(_04540_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10781_ (.A1(_04536_),
    .A2(_04574_),
    .B(_04575_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10782_ (.A1(_04505_),
    .A2(_04534_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10783_ (.A1(_04536_),
    .A2(_04574_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10784_ (.A1(_04505_),
    .A2(_04534_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10785_ (.A1(_04577_),
    .A2(_04578_),
    .B(_04579_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10786_ (.A1(_03830_),
    .A2(_03862_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10787_ (.A1(_04519_),
    .A2(_04532_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10788_ (.A1(_04519_),
    .A2(_04532_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10789_ (.A1(_04521_),
    .A2(_04583_),
    .B(_04584_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10790_ (.A1(_04522_),
    .A2(_04524_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10791_ (.A1(net39),
    .A2(net97),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10792_ (.A1(_04436_),
    .A2(_04587_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10793_ (.A1(_04523_),
    .A2(_04586_),
    .B(_04588_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10794_ (.A1(_04585_),
    .A2(_04589_),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10795_ (.A1(_04581_),
    .A2(_04590_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10796_ (.A1(_04518_),
    .A2(_04533_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10797_ (.A1(_04507_),
    .A2(_04515_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10798_ (.A1(_04529_),
    .A2(_04531_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10799_ (.A1(_04529_),
    .A2(_04531_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10800_ (.A1(_04525_),
    .A2(_04595_),
    .B(_04596_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10801_ (.A1(_04510_),
    .A2(_04514_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10802_ (.A1(net41),
    .A2(net95),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10803_ (.A1(_03871_),
    .A2(net96),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10804_ (.A1(_04587_),
    .A2(_04599_),
    .A3(_04600_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10805_ (.A1(_03907_),
    .A2(_04214_),
    .B1(_04446_),
    .B2(_04235_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10806_ (.A1(_04234_),
    .A2(_03912_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10807_ (.A1(_04530_),
    .A2(_04602_),
    .B1(_04603_),
    .B2(_04447_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10808_ (.A1(_04329_),
    .A2(_04306_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10809_ (.A1(_03902_),
    .A2(_03907_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10810_ (.A1(_04603_),
    .A2(_04606_),
    .A3(_04607_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10811_ (.A1(_04601_),
    .A2(_04605_),
    .A3(_04608_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10812_ (.A1(_04598_),
    .A2(_04609_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10813_ (.A1(_04597_),
    .A2(_04610_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10814_ (.A1(_04190_),
    .A2(_03859_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10815_ (.A1(_03998_),
    .A2(_03945_),
    .B(_04612_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10816_ (.I(net106),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10817_ (.A1(_04614_),
    .A2(_03810_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10818_ (.A1(_04507_),
    .A2(_04616_),
    .Z(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10819_ (.I(_04617_),
    .Z(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10820_ (.A1(_04613_),
    .A2(_04618_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10821_ (.A1(_03866_),
    .A2(_04375_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10822_ (.A1(_03879_),
    .A2(_03958_),
    .B1(_03811_),
    .B2(_03868_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10823_ (.A1(_04363_),
    .A2(_04620_),
    .B1(_04621_),
    .B2(_04511_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10824_ (.A1(_03887_),
    .A2(_04441_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10825_ (.A1(_03877_),
    .A2(_03938_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10826_ (.A1(_04620_),
    .A2(_04623_),
    .A3(_04624_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10827_ (.A1(_04622_),
    .A2(_04625_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10828_ (.A1(_04619_),
    .A2(_04627_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10829_ (.A1(_04594_),
    .A2(_04611_),
    .A3(_04628_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10830_ (.A1(_04592_),
    .A2(_04629_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10831_ (.A1(_04591_),
    .A2(_04630_),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10832_ (.A1(_04576_),
    .A2(_04580_),
    .A3(_04631_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10833_ (.I(_04632_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10834_ (.A1(_04573_),
    .A2(_04633_),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10835_ (.A1(_04570_),
    .A2(_04572_),
    .A3(_04632_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10836_ (.A1(_04634_),
    .A2(_04635_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10837_ (.A1(_04569_),
    .A2(_04636_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10838_ (.A1(_01113_),
    .A2(_04638_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10839_ (.A1(_04555_),
    .A2(_04559_),
    .A3(_04549_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10840_ (.A1(_04555_),
    .A2(_04549_),
    .B(_04559_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10841_ (.A1(_04640_),
    .A2(_04641_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10842_ (.A1(_03863_),
    .A2(_01257_),
    .B1(_00968_),
    .B2(_04470_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10843_ (.I(_04048_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10844_ (.A1(_04644_),
    .A2(_04334_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10845_ (.A1(_04040_),
    .A2(_04552_),
    .A3(_01193_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10846_ (.A1(_04552_),
    .A2(_02822_),
    .B1(_05585_),
    .B2(_04559_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10847_ (.A1(_04643_),
    .A2(_04645_),
    .A3(_04646_),
    .A4(_04647_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10848_ (.A1(_04040_),
    .A2(_01251_),
    .B1(_04642_),
    .B2(_01255_),
    .C(_04649_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10849_ (.A1(_04930_),
    .A2(_04565_),
    .B(_04639_),
    .C(_04650_),
    .ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10850_ (.A1(_03864_),
    .A2(_04562_),
    .B(_04002_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10851_ (.A1(_04003_),
    .A2(_04265_),
    .A3(_04479_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10852_ (.A1(_04087_),
    .A2(_04651_),
    .B(_04652_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10853_ (.A1(_04011_),
    .A2(_04653_),
    .B(_03254_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10854_ (.A1(_04011_),
    .A2(_04653_),
    .B(_04654_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10855_ (.A1(_04545_),
    .A2(_04546_),
    .A3(_04634_),
    .A4(_04635_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10856_ (.A1(_04566_),
    .A2(_04544_),
    .A3(_04635_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10857_ (.A1(_04634_),
    .A2(_04656_),
    .A3(_04657_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10858_ (.A1(_04580_),
    .A2(_04631_),
    .Z(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10859_ (.A1(_04580_),
    .A2(_04631_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10860_ (.A1(_04576_),
    .A2(_04660_),
    .B(_04661_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10861_ (.A1(_03831_),
    .A2(_04041_),
    .A3(_04590_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10862_ (.A1(_04585_),
    .A2(_04589_),
    .B(_04663_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10863_ (.A1(_04592_),
    .A2(_04629_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10864_ (.A1(_04591_),
    .A2(_04630_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10865_ (.A1(_04665_),
    .A2(_04666_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10866_ (.A1(_04096_),
    .A2(_04008_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10867_ (.A1(_04598_),
    .A2(_04609_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10868_ (.A1(_04597_),
    .A2(_04610_),
    .B(_04670_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10869_ (.A1(_04587_),
    .A2(_04600_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10870_ (.A1(net40),
    .A2(net97),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10871_ (.A1(_04524_),
    .A2(_04673_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10872_ (.A1(_04599_),
    .A2(_04672_),
    .B(_04674_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10873_ (.A1(_04671_),
    .A2(_04675_),
    .Z(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10874_ (.A1(_04668_),
    .A2(_04676_),
    .Z(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10875_ (.A1(_04594_),
    .A2(_04628_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(_04594_),
    .A2(_04628_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10877_ (.A1(_04611_),
    .A2(_04678_),
    .B(_04679_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10878_ (.A1(_04613_),
    .A2(_04618_),
    .A3(_04627_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10879_ (.A1(net105),
    .A2(_04375_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10880_ (.A1(_04191_),
    .A2(_04005_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10881_ (.A1(_04616_),
    .A2(_04683_),
    .A3(_04684_),
    .Z(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10882_ (.A1(_03865_),
    .A2(_04307_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10883_ (.A1(_04620_),
    .A2(_04624_),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10884_ (.A1(_04513_),
    .A2(_04686_),
    .B1(_04687_),
    .B2(_04623_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10885_ (.A1(_03886_),
    .A2(_03912_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10886_ (.A1(_04512_),
    .A2(_03920_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10887_ (.A1(_04686_),
    .A2(_04689_),
    .A3(_04690_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10888_ (.A1(_04617_),
    .A2(_04692_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10889_ (.A1(_04685_),
    .A2(_04688_),
    .A3(_04693_),
    .Z(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10890_ (.A1(_04682_),
    .A2(_04694_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10891_ (.A1(_04605_),
    .A2(_04608_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10892_ (.A1(_04605_),
    .A2(_04608_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10893_ (.A1(_04601_),
    .A2(_04696_),
    .B(_04697_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10894_ (.A1(_04622_),
    .A2(_04625_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10895_ (.A1(net42),
    .A2(net95),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10896_ (.I(net41),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10897_ (.A1(_04701_),
    .A2(_03948_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10898_ (.A1(_04673_),
    .A2(_04700_),
    .A3(_04703_),
    .Z(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10899_ (.A1(_03898_),
    .A2(_04433_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10900_ (.A1(_04433_),
    .A2(_04439_),
    .B1(_03913_),
    .B2(_04374_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10901_ (.A1(_04216_),
    .A2(_04705_),
    .B1(_04606_),
    .B2(_04706_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10902_ (.A1(_04393_),
    .A2(_04306_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10903_ (.A1(_03892_),
    .A2(_04439_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10904_ (.A1(_04259_),
    .A2(_04708_),
    .A3(_04709_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10905_ (.A1(_04704_),
    .A2(_04707_),
    .A3(_04710_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10906_ (.A1(_04699_),
    .A2(_04711_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10907_ (.A1(_04698_),
    .A2(_04712_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10908_ (.A1(_04695_),
    .A2(_04714_),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10909_ (.A1(_04681_),
    .A2(_04715_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10910_ (.A1(_04677_),
    .A2(_04716_),
    .Z(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10911_ (.A1(_04667_),
    .A2(_04717_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10912_ (.A1(_04664_),
    .A2(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10913_ (.A1(_04662_),
    .A2(_04719_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10914_ (.A1(_04659_),
    .A2(_04720_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10915_ (.I(_04049_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10916_ (.A1(_04040_),
    .A2(_04041_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10917_ (.A1(_04722_),
    .A2(_04641_),
    .A3(_04723_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10918_ (.A1(_04641_),
    .A2(_04723_),
    .B(_04722_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10919_ (.A1(_04725_),
    .A2(_04726_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10920_ (.I(_03855_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10921_ (.A1(_01792_),
    .A2(_04644_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10922_ (.A1(_04722_),
    .A2(_04729_),
    .B(_04377_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10923_ (.A1(_04728_),
    .A2(_01417_),
    .B1(_05590_),
    .B2(_04552_),
    .C(_04730_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10924_ (.A1(_04006_),
    .A2(_04048_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10925_ (.A1(_04006_),
    .A2(_01493_),
    .B1(_04732_),
    .B2(_01263_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10926_ (.A1(_04644_),
    .A2(_00966_),
    .B(_04731_),
    .C(_04733_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10927_ (.A1(_01430_),
    .A2(_04721_),
    .B1(_04727_),
    .B2(_04097_),
    .C(_04734_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10928_ (.A1(_04655_),
    .A2(_04736_),
    .ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10929_ (.A1(_04662_),
    .A2(_04719_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10930_ (.A1(_04659_),
    .A2(_04720_),
    .B(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10931_ (.A1(_04667_),
    .A2(_04717_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10932_ (.A1(_04664_),
    .A2(_04718_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10933_ (.A1(_03832_),
    .A2(_04009_),
    .A3(_04676_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10934_ (.A1(_04671_),
    .A2(_04675_),
    .B(_04741_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10935_ (.A1(_04681_),
    .A2(_04715_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10936_ (.A1(_04677_),
    .A2(_04716_),
    .B(_04743_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10937_ (.A1(_04096_),
    .A2(_03854_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10938_ (.A1(_04699_),
    .A2(_04711_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10939_ (.A1(_04698_),
    .A2(_04712_),
    .B(_04747_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10940_ (.A1(_04673_),
    .A2(_04703_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10941_ (.A1(_04701_),
    .A2(_04297_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10942_ (.A1(_04600_),
    .A2(_04750_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10943_ (.A1(_04700_),
    .A2(_04749_),
    .B(_04751_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10944_ (.A1(_04748_),
    .A2(_04752_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10945_ (.A1(_04746_),
    .A2(_04753_),
    .Z(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10946_ (.A1(_04613_),
    .A2(_04618_),
    .A3(_04627_),
    .A4(_04694_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10947_ (.A1(_04695_),
    .A2(_04714_),
    .B(_04755_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10948_ (.A1(_04688_),
    .A2(_04693_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10949_ (.A1(_04685_),
    .A2(_04758_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10950_ (.A1(net30),
    .A2(_03851_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10951_ (.A1(net107),
    .A2(_03809_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10952_ (.A1(net105),
    .A2(net33),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10953_ (.A1(net106),
    .A2(_03956_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10954_ (.A1(_04761_),
    .A2(_04762_),
    .A3(_04763_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10955_ (.A1(_04760_),
    .A2(_04764_),
    .Z(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10956_ (.A1(_04686_),
    .A2(_04690_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10957_ (.A1(_03865_),
    .A2(net34),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10958_ (.A1(_04624_),
    .A2(_04768_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10959_ (.A1(_04689_),
    .A2(_04766_),
    .B(_04769_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10960_ (.A1(_04190_),
    .A2(_04004_),
    .B1(_03859_),
    .B2(_04231_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10961_ (.A1(_04612_),
    .A2(_04761_),
    .B1(_04771_),
    .B2(_04683_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10962_ (.A1(net101),
    .A2(_04257_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10963_ (.A1(_04512_),
    .A2(_04214_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10964_ (.A1(_04768_),
    .A2(_04773_),
    .A3(_04774_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10965_ (.A1(_04772_),
    .A2(_04775_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10966_ (.A1(_04770_),
    .A2(_04776_),
    .Z(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10967_ (.A1(_04765_),
    .A2(_04777_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10968_ (.I(_04704_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10969_ (.A1(_04707_),
    .A2(_04710_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10970_ (.A1(_04707_),
    .A2(_04710_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10971_ (.A1(_04780_),
    .A2(_04781_),
    .B(_04782_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10972_ (.A1(_04618_),
    .A2(_04692_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10973_ (.A1(_04617_),
    .A2(_04692_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10974_ (.A1(_04688_),
    .A2(_04784_),
    .B(_04785_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10975_ (.A1(_04007_),
    .A2(_03841_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10976_ (.A1(net42),
    .A2(_03948_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10977_ (.A1(_04750_),
    .A2(_04788_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10978_ (.A1(_04787_),
    .A2(_04790_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10979_ (.A1(_03898_),
    .A2(_04433_),
    .B1(_03908_),
    .B2(_03892_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10980_ (.A1(_04329_),
    .A2(_04234_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10981_ (.A1(_04708_),
    .A2(_04792_),
    .B1(_04793_),
    .B2(_04607_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10982_ (.A1(net40),
    .A2(net98),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10983_ (.A1(_04393_),
    .A2(_03907_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10984_ (.A1(_04793_),
    .A2(_04795_),
    .A3(_04796_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10985_ (.A1(_04794_),
    .A2(_04797_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10986_ (.A1(_04791_),
    .A2(_04798_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10987_ (.A1(_04783_),
    .A2(_04786_),
    .A3(_04799_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10988_ (.A1(_04759_),
    .A2(_04779_),
    .A3(_04801_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10989_ (.A1(_04757_),
    .A2(_04802_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10990_ (.A1(_04754_),
    .A2(_04803_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10991_ (.A1(_04744_),
    .A2(_04804_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10992_ (.A1(_04742_),
    .A2(_04805_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10993_ (.A1(_04739_),
    .A2(_04740_),
    .B(_04806_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10994_ (.A1(_04739_),
    .A2(_04740_),
    .A3(_04806_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10995_ (.A1(_04807_),
    .A2(_04808_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10996_ (.A1(_04738_),
    .A2(_04809_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10997_ (.A1(_04732_),
    .A2(_04726_),
    .B(_04039_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10998_ (.I(_04039_),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10999_ (.A1(_04732_),
    .A2(_04813_),
    .A3(_04726_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11000_ (.A1(_04812_),
    .A2(_04814_),
    .Z(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11001_ (.I(_04020_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11002_ (.I(_04816_),
    .Z(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11003_ (.A1(_03853_),
    .A2(_04728_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11004_ (.I(_04818_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11005_ (.A1(_04817_),
    .A2(_04637_),
    .B1(_02692_),
    .B2(_04819_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11006_ (.A1(_03857_),
    .A2(_01418_),
    .B1(_01410_),
    .B2(_04644_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11007_ (.A1(_04728_),
    .A2(_05517_),
    .B1(_05520_),
    .B2(_04813_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11008_ (.A1(_04820_),
    .A2(_04821_),
    .A3(_04823_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11009_ (.A1(_03853_),
    .A2(_05498_),
    .B1(_04815_),
    .B2(_05503_),
    .C(_04824_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11010_ (.A1(_04012_),
    .A2(_04048_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11011_ (.A1(_04722_),
    .A2(_04651_),
    .B(_04826_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11012_ (.A1(_04265_),
    .A2(_04479_),
    .B(_04827_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11013_ (.A1(_04014_),
    .A2(_04055_),
    .B(_04828_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11014_ (.A1(_04813_),
    .A2(_04829_),
    .B(_04271_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11015_ (.A1(_04813_),
    .A2(_04829_),
    .B(_04830_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11016_ (.A1(_00675_),
    .A2(_04810_),
    .B(_04825_),
    .C(_04831_),
    .ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11017_ (.A1(_04023_),
    .A2(_04816_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11018_ (.I(_04833_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11019_ (.A1(_04015_),
    .A2(_04827_),
    .B(_03858_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11020_ (.A1(_04027_),
    .A2(_04051_),
    .B(_04835_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11021_ (.A1(_04016_),
    .A2(_04108_),
    .B(_04836_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11022_ (.A1(_04834_),
    .A2(_04837_),
    .B(_01488_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11023_ (.A1(_04834_),
    .A2(_04837_),
    .B(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11024_ (.A1(_04018_),
    .A2(_04816_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11025_ (.A1(_04018_),
    .A2(_04171_),
    .B1(_04840_),
    .B2(_04215_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11026_ (.I(_03847_),
    .Z(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11027_ (.A1(_01792_),
    .A2(_04817_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11028_ (.A1(_04834_),
    .A2(_04844_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11029_ (.A1(_03857_),
    .A2(_01858_),
    .A3(_04065_),
    .B1(_04626_),
    .B2(_04817_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11030_ (.A1(_04842_),
    .A2(_00233_),
    .B1(_04845_),
    .B2(_04604_),
    .C(_04846_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11031_ (.A1(_04659_),
    .A2(_04720_),
    .A3(_04809_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11032_ (.A1(_04739_),
    .A2(_04740_),
    .A3(_04806_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11033_ (.A1(_04737_),
    .A2(_04807_),
    .B(_04849_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11034_ (.A1(_04744_),
    .A2(_04804_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11035_ (.A1(_04742_),
    .A2(_04805_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11036_ (.A1(_04851_),
    .A2(_04852_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11037_ (.A1(_03831_),
    .A2(_03855_),
    .A3(_04753_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11038_ (.A1(_04748_),
    .A2(_04752_),
    .B(_04855_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11039_ (.A1(_04757_),
    .A2(_04802_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11040_ (.A1(_04754_),
    .A2(_04803_),
    .B(_04857_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11041_ (.A1(_04786_),
    .A2(_04799_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11042_ (.A1(_04786_),
    .A2(_04799_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11043_ (.A1(_04783_),
    .A2(_04859_),
    .B(_04860_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11044_ (.A1(_03861_),
    .A2(_04297_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11045_ (.A1(_04703_),
    .A2(_04862_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11046_ (.A1(_04787_),
    .A2(_04790_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11047_ (.A1(_04863_),
    .A2(_04864_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11048_ (.A1(_04861_),
    .A2(_04866_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11049_ (.A1(_04096_),
    .A2(_04019_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11050_ (.A1(_04867_),
    .A2(_04868_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11051_ (.A1(_04759_),
    .A2(_04779_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11052_ (.I(_04801_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11053_ (.A1(_04759_),
    .A2(_04779_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11054_ (.A1(_04870_),
    .A2(_04871_),
    .B(_04872_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11055_ (.A1(_04794_),
    .A2(_04797_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11056_ (.A1(_04791_),
    .A2(_04798_),
    .B(_04874_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11057_ (.A1(_04772_),
    .A2(_04775_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11058_ (.A1(_04770_),
    .A2(_04776_),
    .B(_04877_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11059_ (.A1(_03854_),
    .A2(_04295_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11060_ (.A1(net43),
    .A2(_03948_),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11061_ (.A1(_04862_),
    .A2(_04880_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11062_ (.A1(_04879_),
    .A2(_04881_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11063_ (.A1(_04393_),
    .A2(_04235_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11064_ (.A1(_04793_),
    .A2(_04796_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11065_ (.A1(_04709_),
    .A2(_04883_),
    .B1(_04884_),
    .B2(_04795_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11066_ (.A1(_04701_),
    .A2(_04306_),
    .Z(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11067_ (.A1(_03872_),
    .A2(_04439_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11068_ (.A1(_04883_),
    .A2(_04886_),
    .A3(_04888_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11069_ (.A1(_04885_),
    .A2(_04889_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11070_ (.A1(_04882_),
    .A2(_04890_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11071_ (.A1(_04875_),
    .A2(_04878_),
    .A3(_04891_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11072_ (.A1(_04765_),
    .A2(_04777_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11073_ (.A1(_04760_),
    .A2(_04764_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11074_ (.A1(_04190_),
    .A2(_04017_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11075_ (.A1(_03851_),
    .A2(_04231_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11076_ (.A1(net109),
    .A2(net31),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11077_ (.A1(_04760_),
    .A2(_04897_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11078_ (.A1(_04895_),
    .A2(_04896_),
    .B(_04899_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11079_ (.A1(_03987_),
    .A2(_04441_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11080_ (.A1(net107),
    .A2(net32),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11081_ (.A1(net106),
    .A2(_03937_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11082_ (.A1(_04902_),
    .A2(_04903_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11083_ (.A1(_04901_),
    .A2(_04904_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11084_ (.A1(_04894_),
    .A2(_04900_),
    .A3(_04905_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11085_ (.A1(_04768_),
    .A2(_04774_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11086_ (.A1(net104),
    .A2(net35),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11087_ (.A1(_04690_),
    .A2(_04908_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11088_ (.A1(_04773_),
    .A2(_04907_),
    .B(_04909_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11089_ (.A1(_04614_),
    .A2(_04309_),
    .B1(_03810_),
    .B2(_04004_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11090_ (.A1(_04616_),
    .A2(_04902_),
    .B1(_04911_),
    .B2(_04762_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11091_ (.A1(_04512_),
    .A2(_03902_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11092_ (.A1(_04330_),
    .A2(_04908_),
    .A3(_04913_),
    .Z(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11093_ (.A1(_04912_),
    .A2(_04914_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11094_ (.A1(_04910_),
    .A2(_04915_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11095_ (.A1(_04906_),
    .A2(_04916_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11096_ (.A1(_04893_),
    .A2(_04917_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11097_ (.A1(_04892_),
    .A2(_04918_),
    .Z(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11098_ (.A1(_04873_),
    .A2(_04920_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11099_ (.A1(_04869_),
    .A2(_04921_),
    .Z(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11100_ (.A1(_04858_),
    .A2(_04922_),
    .Z(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11101_ (.A1(_04856_),
    .A2(_04923_),
    .Z(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11102_ (.A1(_04853_),
    .A2(_04924_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11103_ (.A1(_04848_),
    .A2(_04850_),
    .A3(_04925_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11104_ (.A1(_04848_),
    .A2(_04850_),
    .B(_04925_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11105_ (.A1(_00992_),
    .A2(_04927_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11106_ (.A1(_04812_),
    .A2(_04818_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11107_ (.A1(_04834_),
    .A2(_04929_),
    .Z(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11108_ (.A1(_05431_),
    .A2(_04931_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11109_ (.A1(_04926_),
    .A2(_04928_),
    .B(_04932_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11110_ (.A1(_04839_),
    .A2(_04841_),
    .A3(_04847_),
    .A4(_04933_),
    .ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11111_ (.A1(_04853_),
    .A2(_04924_),
    .Z(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11112_ (.A1(_04934_),
    .A2(_04927_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11113_ (.A1(_03831_),
    .A2(_04019_),
    .A3(_04867_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11114_ (.A1(_04861_),
    .A2(_04866_),
    .B(_04936_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11115_ (.A1(_04873_),
    .A2(_04920_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11116_ (.A1(_04869_),
    .A2(_04921_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11117_ (.A1(_04938_),
    .A2(_04939_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11118_ (.A1(_04878_),
    .A2(_04891_),
    .Z(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11119_ (.A1(_04878_),
    .A2(_04891_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11120_ (.A1(_04875_),
    .A2(_04942_),
    .B(_04943_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11121_ (.A1(_04862_),
    .A2(_04880_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11122_ (.A1(_04879_),
    .A2(_04881_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11123_ (.A1(_04945_),
    .A2(_04946_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11124_ (.A1(_04944_),
    .A2(_04947_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11125_ (.A1(_03830_),
    .A2(_03847_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11126_ (.A1(_04948_),
    .A2(_04949_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11127_ (.A1(_04893_),
    .A2(_04917_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11128_ (.A1(_04892_),
    .A2(_04918_),
    .B(_04952_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11129_ (.A1(_04885_),
    .A2(_04889_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11130_ (.A1(_04882_),
    .A2(_04890_),
    .B(_04954_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11131_ (.A1(_04332_),
    .A2(_04908_),
    .A3(_04913_),
    .Z(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11132_ (.A1(_04912_),
    .A2(_04956_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11133_ (.A1(_04910_),
    .A2(_04915_),
    .B(_04957_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11134_ (.A1(net45),
    .A2(_04295_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11135_ (.A1(net44),
    .A2(_04183_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11136_ (.A1(_04880_),
    .A2(_04960_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11137_ (.A1(_04008_),
    .A2(_03932_),
    .B1(_04123_),
    .B2(net44),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11138_ (.A1(_04961_),
    .A2(_04963_),
    .Z(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11139_ (.A1(_04959_),
    .A2(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11140_ (.A1(_04883_),
    .A2(_04888_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11141_ (.A1(_03871_),
    .A2(_04235_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11142_ (.A1(_04796_),
    .A2(_04967_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11143_ (.A1(_04886_),
    .A2(_04966_),
    .B(_04968_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11144_ (.A1(_03861_),
    .A2(_03923_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11145_ (.A1(_04701_),
    .A2(_04194_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11146_ (.A1(_04967_),
    .A2(_04971_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11147_ (.A1(_04970_),
    .A2(_04972_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11148_ (.A1(_04969_),
    .A2(_04974_),
    .Z(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11149_ (.A1(_04969_),
    .A2(_04974_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11150_ (.A1(_04975_),
    .A2(_04976_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11151_ (.A1(_04965_),
    .A2(_04977_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11152_ (.A1(_04955_),
    .A2(_04958_),
    .A3(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11153_ (.A1(_04900_),
    .A2(_04905_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11154_ (.A1(_04900_),
    .A2(_04905_),
    .Z(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11155_ (.A1(_04894_),
    .A2(_04980_),
    .A3(_04981_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11156_ (.A1(_04906_),
    .A2(_04916_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11157_ (.A1(_04982_),
    .A2(_04983_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11158_ (.A1(net108),
    .A2(net32),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11159_ (.A1(net30),
    .A2(net110),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11160_ (.A1(_04897_),
    .A2(_04986_),
    .A3(_04987_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11161_ (.A1(_04899_),
    .A2(_04988_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11162_ (.A1(net107),
    .A2(_03937_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11163_ (.A1(net105),
    .A2(net35),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11164_ (.A1(_04614_),
    .A2(_04446_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11165_ (.A1(_04990_),
    .A2(_04991_),
    .A3(_04992_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11166_ (.A1(_04989_),
    .A2(_04993_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11167_ (.A1(_04980_),
    .A2(_04994_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11168_ (.A1(net104),
    .A2(_04257_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11169_ (.A1(_04908_),
    .A2(_04913_),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11170_ (.A1(_04774_),
    .A2(_04997_),
    .B1(_04998_),
    .B2(_04331_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11171_ (.A1(_04763_),
    .A2(_04990_),
    .B1(_04904_),
    .B2(_04901_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11172_ (.A1(_03882_),
    .A2(_03887_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11173_ (.A1(net103),
    .A2(net37),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11174_ (.A1(_04997_),
    .A2(_05002_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11175_ (.A1(_05001_),
    .A2(_05003_),
    .Z(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11176_ (.A1(_05000_),
    .A2(_05004_),
    .Z(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11177_ (.A1(_04999_),
    .A2(_05005_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11178_ (.A1(_04996_),
    .A2(_05007_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11179_ (.A1(_04985_),
    .A2(_05008_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11180_ (.A1(_04979_),
    .A2(_05009_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11181_ (.A1(_04953_),
    .A2(_05010_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11182_ (.A1(_04950_),
    .A2(_05011_),
    .Z(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11183_ (.A1(_04937_),
    .A2(_04941_),
    .A3(_05012_),
    .Z(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11184_ (.A1(_04858_),
    .A2(_04922_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11185_ (.A1(_04856_),
    .A2(_04923_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11186_ (.A1(_05014_),
    .A2(_05015_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11187_ (.A1(_05013_),
    .A2(_05016_),
    .Z(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11188_ (.A1(_04935_),
    .A2(_05018_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11189_ (.A1(_04935_),
    .A2(_05018_),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11190_ (.A1(_01113_),
    .A2(_05020_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11191_ (.I(_03850_),
    .Z(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11192_ (.A1(_04022_),
    .A2(_04929_),
    .B(_04840_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11193_ (.A1(_05022_),
    .A2(_05023_),
    .B(_00045_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11194_ (.A1(_05022_),
    .A2(_05023_),
    .B(_05024_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11195_ (.I(_03849_),
    .Z(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11196_ (.A1(_04023_),
    .A2(_04816_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11197_ (.A1(_04833_),
    .A2(_04835_),
    .B(_05027_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11198_ (.A1(_05022_),
    .A2(_05029_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11199_ (.A1(_04026_),
    .A2(_04025_),
    .B1(_04055_),
    .B2(_05030_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11200_ (.A1(_04756_),
    .A2(_05031_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11201_ (.A1(_04842_),
    .A2(_05026_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11202_ (.A1(_03848_),
    .A2(_01418_),
    .B1(_05507_),
    .B2(_04817_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11203_ (.A1(_05202_),
    .A2(_03847_),
    .A3(_05026_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11204_ (.A1(_04842_),
    .A2(_05026_),
    .B(_04593_),
    .C(_05035_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11205_ (.A1(_00959_),
    .A2(_05033_),
    .B(_05034_),
    .C(_05036_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11206_ (.A1(_05026_),
    .A2(_04171_),
    .B(_05032_),
    .C(_05037_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11207_ (.A1(_05019_),
    .A2(_05021_),
    .B(_05025_),
    .C(_05038_),
    .ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11208_ (.A1(_04944_),
    .A2(_04947_),
    .Z(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11209_ (.A1(_04948_),
    .A2(_04949_),
    .B(_05040_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11210_ (.A1(_04953_),
    .A2(_05010_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11211_ (.I(_05011_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11212_ (.A1(_04950_),
    .A2(_05043_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11213_ (.A1(_05042_),
    .A2(_05044_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11214_ (.A1(_04958_),
    .A2(_04978_),
    .Z(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11215_ (.A1(_04958_),
    .A2(_04978_),
    .Z(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11216_ (.A1(_04955_),
    .A2(_05046_),
    .B(_05047_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11217_ (.A1(_04959_),
    .A2(_04964_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11218_ (.A1(_04961_),
    .A2(_05050_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11219_ (.A1(_05048_),
    .A2(_05051_),
    .Z(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11220_ (.A1(_04985_),
    .A2(_05008_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11221_ (.A1(_04979_),
    .A2(_05009_),
    .B(_05053_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11222_ (.A1(_04980_),
    .A2(_04994_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11223_ (.A1(_04996_),
    .A2(_05007_),
    .B(_05055_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11224_ (.A1(_04899_),
    .A2(_04988_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11225_ (.A1(_04989_),
    .A2(_04993_),
    .B(_05057_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11226_ (.A1(net110),
    .A2(net31),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11227_ (.A1(_04897_),
    .A2(_04987_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11228_ (.A1(_04895_),
    .A2(_05059_),
    .B1(_05061_),
    .B2(_04986_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11229_ (.A1(_03851_),
    .A2(_04307_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11230_ (.A1(net109),
    .A2(net32),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11231_ (.A1(_05059_),
    .A2(_05064_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11232_ (.A1(_05063_),
    .A2(_05065_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11233_ (.A1(_05062_),
    .A2(_05066_),
    .Z(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11234_ (.A1(_03987_),
    .A2(_03903_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11235_ (.A1(_04004_),
    .A2(_04446_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11236_ (.A1(_04614_),
    .A2(_04214_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11237_ (.A1(_05069_),
    .A2(_05070_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11238_ (.A1(_05068_),
    .A2(_05072_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11239_ (.A1(_05067_),
    .A2(_05073_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11240_ (.A1(_05058_),
    .A2(_05074_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11241_ (.A1(_03866_),
    .A2(_04329_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11242_ (.A1(_04913_),
    .A2(_05076_),
    .B1(_05003_),
    .B2(_05001_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11243_ (.I(_05077_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11244_ (.A1(_04990_),
    .A2(_04992_),
    .Z(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11245_ (.A1(_04903_),
    .A2(_05069_),
    .B1(_05079_),
    .B2(_04991_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11246_ (.A1(_04394_),
    .A2(_05076_),
    .Z(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11247_ (.A1(_03872_),
    .A2(_03888_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11248_ (.A1(_05081_),
    .A2(_05083_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11249_ (.A1(_05080_),
    .A2(_05084_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11250_ (.A1(_05078_),
    .A2(_05085_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11251_ (.A1(_05075_),
    .A2(_05086_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11252_ (.A1(_05056_),
    .A2(_05087_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11253_ (.A1(_04965_),
    .A2(_04977_),
    .B(_04975_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11254_ (.A1(_05000_),
    .A2(_05004_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11255_ (.A1(_04999_),
    .A2(_05005_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11256_ (.A1(_05090_),
    .A2(_05091_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11257_ (.A1(net46),
    .A2(_03842_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11258_ (.A1(net45),
    .A2(_03950_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11259_ (.A1(_04960_),
    .A2(_05095_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11260_ (.A1(_05094_),
    .A2(_05096_),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11261_ (.A1(_03991_),
    .A2(_04374_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11262_ (.A1(_04888_),
    .A2(_05098_),
    .B1(_04972_),
    .B2(_04970_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11263_ (.A1(_04007_),
    .A2(_03923_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11264_ (.A1(net42),
    .A2(_04194_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11265_ (.A1(_05098_),
    .A2(_05101_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11266_ (.A1(_05100_),
    .A2(_05102_),
    .Z(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11267_ (.A1(_05099_),
    .A2(_05103_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11268_ (.A1(_05097_),
    .A2(_05105_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11269_ (.A1(_05092_),
    .A2(_05106_),
    .Z(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11270_ (.A1(_05089_),
    .A2(_05107_),
    .Z(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11271_ (.A1(_05088_),
    .A2(_05108_),
    .Z(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11272_ (.A1(_05054_),
    .A2(_05109_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11273_ (.A1(_05052_),
    .A2(_05110_),
    .Z(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11274_ (.A1(_05041_),
    .A2(_05045_),
    .A3(_05111_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11275_ (.I(_04941_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11276_ (.A1(_05113_),
    .A2(_05012_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11277_ (.A1(_05113_),
    .A2(_05012_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11278_ (.A1(_04937_),
    .A2(_05114_),
    .B(_05116_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11279_ (.A1(_05112_),
    .A2(_05117_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11280_ (.A1(_05014_),
    .A2(_05015_),
    .B(_05013_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11281_ (.A1(_05014_),
    .A2(_05015_),
    .A3(_05013_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11282_ (.A1(_04934_),
    .A2(_05119_),
    .B(_05120_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11283_ (.A1(_04850_),
    .A2(_05121_),
    .Z(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11284_ (.A1(_04925_),
    .A2(_05018_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11285_ (.A1(_04848_),
    .A2(_05122_),
    .B1(_05123_),
    .B2(_05121_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11286_ (.A1(_05118_),
    .A2(_05124_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11287_ (.A1(_05022_),
    .A2(_05023_),
    .B(_05033_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11288_ (.A1(_04842_),
    .A2(_00585_),
    .B1(_05127_),
    .B2(_01255_),
    .C(_00588_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11289_ (.A1(_05115_),
    .A2(_05125_),
    .B(_05128_),
    .ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11290_ (.A1(_05112_),
    .A2(_05117_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11291_ (.A1(_04848_),
    .A2(_05122_),
    .B1(_05123_),
    .B2(_05121_),
    .C(_05118_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11292_ (.A1(_05129_),
    .A2(_05130_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11293_ (.A1(_05048_),
    .A2(_05051_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11294_ (.A1(_05054_),
    .A2(_05109_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11295_ (.A1(_05052_),
    .A2(_05110_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11296_ (.A1(_05133_),
    .A2(_05134_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11297_ (.I(_05106_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11298_ (.I(_05089_),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11299_ (.A1(_05138_),
    .A2(_05107_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11300_ (.A1(_05092_),
    .A2(_05137_),
    .B(_05139_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11301_ (.A1(_04960_),
    .A2(_05095_),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11302_ (.A1(_05094_),
    .A2(_05096_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11303_ (.A1(_05141_),
    .A2(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11304_ (.A1(_05140_),
    .A2(_05143_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11305_ (.A1(_05056_),
    .A2(_05087_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11306_ (.A1(_05088_),
    .A2(_05108_),
    .B(_05145_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11307_ (.A1(_05058_),
    .A2(_05074_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11308_ (.A1(_05075_),
    .A2(_05086_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11309_ (.A1(_05148_),
    .A2(_05149_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11310_ (.A1(_05062_),
    .A2(_05066_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11311_ (.A1(_05067_),
    .A2(_05073_),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11312_ (.A1(_05151_),
    .A2(_05152_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11313_ (.A1(net110),
    .A2(_04309_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11314_ (.A1(_04897_),
    .A2(_05154_),
    .B1(_05065_),
    .B2(_05063_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11315_ (.A1(_03852_),
    .A2(_03926_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11316_ (.A1(_04017_),
    .A2(_03938_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11317_ (.A1(_05154_),
    .A2(_05157_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11318_ (.A1(_05156_),
    .A2(_05159_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11319_ (.A1(_05155_),
    .A2(_05160_),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11320_ (.A1(_04005_),
    .A2(_03914_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11321_ (.A1(_03989_),
    .A2(_03893_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11322_ (.A1(_03859_),
    .A2(_03904_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11323_ (.A1(_05162_),
    .A2(_05163_),
    .A3(_05164_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11324_ (.A1(_05161_),
    .A2(_05165_),
    .Z(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11325_ (.A1(_05153_),
    .A2(_05166_),
    .Z(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11326_ (.A1(_03868_),
    .A2(_03883_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11327_ (.A1(_05002_),
    .A2(_05168_),
    .B1(_05081_),
    .B2(_05083_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11328_ (.A1(_05069_),
    .A2(_05070_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11329_ (.A1(_05068_),
    .A2(_05072_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11330_ (.A1(_05171_),
    .A2(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11331_ (.A1(_03991_),
    .A2(_03888_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11332_ (.A1(_03872_),
    .A2(_03879_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11333_ (.A1(_05168_),
    .A2(_05175_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11334_ (.A1(_05174_),
    .A2(_05176_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11335_ (.A1(_05173_),
    .A2(_05177_),
    .Z(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11336_ (.A1(_05170_),
    .A2(_05178_),
    .Z(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11337_ (.A1(_05167_),
    .A2(_05179_),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11338_ (.A1(_05099_),
    .A2(_05103_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11339_ (.A1(_05097_),
    .A2(_05105_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11340_ (.A1(_05182_),
    .A2(_05183_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11341_ (.A1(_05080_),
    .A2(_05084_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11342_ (.A1(_05078_),
    .A2(_05085_),
    .B(_05185_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11343_ (.A1(_04019_),
    .A2(_03934_),
    .B1(_03952_),
    .B2(net46),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11344_ (.A1(net46),
    .A2(_03934_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11345_ (.A1(_05095_),
    .A2(_05188_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11346_ (.A1(_05187_),
    .A2(_05189_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11347_ (.A1(_03861_),
    .A2(_04237_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11348_ (.A1(_04971_),
    .A2(_05192_),
    .B1(_05102_),
    .B2(_05100_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11349_ (.A1(_03854_),
    .A2(_03924_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11350_ (.A1(_04007_),
    .A2(_04195_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11351_ (.A1(_05192_),
    .A2(_05195_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11352_ (.A1(_05194_),
    .A2(_05196_),
    .Z(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11353_ (.A1(_05193_),
    .A2(_05197_),
    .Z(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11354_ (.A1(_05190_),
    .A2(_05198_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11355_ (.A1(_05186_),
    .A2(_05199_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11356_ (.A1(_05184_),
    .A2(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11357_ (.A1(_05150_),
    .A2(_05181_),
    .A3(_05201_),
    .Z(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11358_ (.A1(_05146_),
    .A2(_05203_),
    .Z(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11359_ (.A1(_05144_),
    .A2(_05204_),
    .Z(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11360_ (.A1(_05132_),
    .A2(_05135_),
    .A3(_05205_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11361_ (.A1(_05045_),
    .A2(_05111_),
    .Z(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11362_ (.A1(_05045_),
    .A2(_05111_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11363_ (.A1(_05041_),
    .A2(_05207_),
    .B(_05208_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11364_ (.A1(_05206_),
    .A2(_05209_),
    .Z(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11365_ (.A1(_05131_),
    .A2(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11366_ (.A1(_05131_),
    .A2(_05210_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11367_ (.A1(_00671_),
    .A2(_05212_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11368_ (.A1(_05211_),
    .A2(_05214_),
    .B(_00674_),
    .ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11369_ (.I(_05209_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11370_ (.A1(_05206_),
    .A2(_05215_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11371_ (.A1(_05131_),
    .A2(_05210_),
    .B(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11372_ (.A1(_05133_),
    .A2(_05134_),
    .A3(_05205_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11373_ (.A1(_05133_),
    .A2(_05134_),
    .B(_05205_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11374_ (.A1(_05132_),
    .A2(_05218_),
    .B(_05219_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11375_ (.I(_05144_),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11376_ (.I(_05203_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11377_ (.A1(_05146_),
    .A2(_05222_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11378_ (.A1(_05221_),
    .A2(_05204_),
    .B(_05224_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11379_ (.A1(_05170_),
    .A2(_05178_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11380_ (.A1(_05173_),
    .A2(_05177_),
    .B(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11381_ (.A1(_04008_),
    .A2(_03899_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11382_ (.A1(_05101_),
    .A2(_05228_),
    .B1(_05196_),
    .B2(_05194_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11383_ (.A1(_04020_),
    .A2(_03975_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11384_ (.A1(_05188_),
    .A2(_05228_),
    .A3(_05230_),
    .Z(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11385_ (.A1(_05227_),
    .A2(_05229_),
    .A3(_05231_),
    .Z(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11386_ (.A1(_05225_),
    .A2(_05232_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11387_ (.A1(_05193_),
    .A2(_05197_),
    .B1(_05198_),
    .B2(_05190_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11388_ (.A1(_04728_),
    .A2(_03910_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11389_ (.A1(_05150_),
    .A2(_05181_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11390_ (.A1(_05150_),
    .A2(_05181_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11391_ (.A1(_05237_),
    .A2(_05201_),
    .B(_05238_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11392_ (.A1(_05186_),
    .A2(_05199_),
    .Z(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11393_ (.A1(_05184_),
    .A2(_05200_),
    .B(_05240_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11394_ (.A1(_05189_),
    .A2(_05241_),
    .Z(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11395_ (.A1(_05140_),
    .A2(_05143_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11396_ (.A1(_05153_),
    .A2(_05166_),
    .Z(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11397_ (.A1(_05167_),
    .A2(_05179_),
    .B(_05244_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11398_ (.I(_05160_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11399_ (.A1(_05155_),
    .A2(_05247_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11400_ (.A1(_05161_),
    .A2(_05165_),
    .B(_05248_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11401_ (.A1(_03849_),
    .A2(_03941_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11402_ (.A1(_03989_),
    .A2(_03883_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11403_ (.A1(_03862_),
    .A2(_03890_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11404_ (.A1(_05250_),
    .A2(_05251_),
    .A3(_05252_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11405_ (.A1(_05249_),
    .A2(_05253_),
    .Z(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11406_ (.A1(_04394_),
    .A2(_04471_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11407_ (.A1(_03992_),
    .A2(_03890_),
    .A3(_05176_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11408_ (.I0(_04472_),
    .I1(_05255_),
    .S(_05257_),
    .Z(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11409_ (.A1(_03852_),
    .A2(_03915_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11410_ (.A1(_04017_),
    .A2(_03928_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11411_ (.A1(_03860_),
    .A2(_03894_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11412_ (.A1(_05064_),
    .A2(_05250_),
    .B1(_05159_),
    .B2(_05156_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11413_ (.A1(_05260_),
    .A2(_05261_),
    .A3(_05262_),
    .Z(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11414_ (.A1(_04005_),
    .A2(_03904_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11415_ (.A1(_05162_),
    .A2(_05164_),
    .Z(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11416_ (.A1(_05070_),
    .A2(_05264_),
    .B1(_05265_),
    .B2(_05163_),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11417_ (.A1(_03992_),
    .A2(_03880_),
    .ZN(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11418_ (.A1(_05264_),
    .A2(_05266_),
    .A3(_05268_),
    .Z(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11419_ (.A1(_05259_),
    .A2(_05263_),
    .A3(_05269_),
    .Z(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11420_ (.A1(_05254_),
    .A2(_05258_),
    .A3(_05270_),
    .Z(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11421_ (.A1(_05243_),
    .A2(_05246_),
    .A3(_05271_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11422_ (.A1(_05239_),
    .A2(_05242_),
    .A3(_05272_),
    .Z(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11423_ (.A1(_05235_),
    .A2(_05236_),
    .A3(_05273_),
    .Z(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11424_ (.A1(_05220_),
    .A2(_05233_),
    .A3(_05274_),
    .Z(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11425_ (.A1(_05217_),
    .A2(_05275_),
    .Z(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11426_ (.A1(_05217_),
    .A2(_05275_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11427_ (.A1(_02152_),
    .A2(_05276_),
    .A3(_05277_),
    .B(_00735_),
    .ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(Operation[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(Operation[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(Operation[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(Operation[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(a_operand[0]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(a_operand[10]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(a_operand[11]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(a_operand[12]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input9 (.I(a_operand[13]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(a_operand[14]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input11 (.I(a_operand[15]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input12 (.I(a_operand[16]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input13 (.I(a_operand[17]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(a_operand[18]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(a_operand[19]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(a_operand[1]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input17 (.I(a_operand[20]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(a_operand[21]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input19 (.I(a_operand[22]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(a_operand[23]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input21 (.I(a_operand[24]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input22 (.I(a_operand[25]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input23 (.I(a_operand[26]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input24 (.I(a_operand[27]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(a_operand[28]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input26 (.I(a_operand[29]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input27 (.I(a_operand[2]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input28 (.I(a_operand[30]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input29 (.I(a_operand[31]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input30 (.I(a_operand[32]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input31 (.I(a_operand[33]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(a_operand[34]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input33 (.I(a_operand[35]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input34 (.I(a_operand[36]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input35 (.I(a_operand[37]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input36 (.I(a_operand[38]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input37 (.I(a_operand[39]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input38 (.I(a_operand[3]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input39 (.I(a_operand[40]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(a_operand[41]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input41 (.I(a_operand[42]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(a_operand[43]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input43 (.I(a_operand[44]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input44 (.I(a_operand[45]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input45 (.I(a_operand[46]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(a_operand[47]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input47 (.I(a_operand[48]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input48 (.I(a_operand[49]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(a_operand[4]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input50 (.I(a_operand[50]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input51 (.I(a_operand[51]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(a_operand[52]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input53 (.I(a_operand[53]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input54 (.I(a_operand[54]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input55 (.I(a_operand[55]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(a_operand[56]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input57 (.I(a_operand[57]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input58 (.I(a_operand[58]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input59 (.I(a_operand[59]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input60 (.I(a_operand[5]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input61 (.I(a_operand[60]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input62 (.I(a_operand[61]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input63 (.I(a_operand[62]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input64 (.I(a_operand[63]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input65 (.I(a_operand[6]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(a_operand[7]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input67 (.I(a_operand[8]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input68 (.I(a_operand[9]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(b_operand[0]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input70 (.I(b_operand[10]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(b_operand[11]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input72 (.I(b_operand[12]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input73 (.I(b_operand[13]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input74 (.I(b_operand[14]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input75 (.I(b_operand[15]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input76 (.I(b_operand[16]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(b_operand[17]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(b_operand[18]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input79 (.I(b_operand[19]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input80 (.I(b_operand[1]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(b_operand[20]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input82 (.I(b_operand[21]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input83 (.I(b_operand[22]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input84 (.I(b_operand[23]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input85 (.I(b_operand[24]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input86 (.I(b_operand[25]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input87 (.I(b_operand[26]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input88 (.I(b_operand[27]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input89 (.I(b_operand[28]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input90 (.I(b_operand[29]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input91 (.I(b_operand[2]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input92 (.I(b_operand[30]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input93 (.I(b_operand[31]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input94 (.I(b_operand[32]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input95 (.I(b_operand[33]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input96 (.I(b_operand[34]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input97 (.I(b_operand[35]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input98 (.I(b_operand[36]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input99 (.I(b_operand[37]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input100 (.I(b_operand[38]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input101 (.I(b_operand[39]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input102 (.I(b_operand[3]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input103 (.I(b_operand[40]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input104 (.I(b_operand[41]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input105 (.I(b_operand[42]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input106 (.I(b_operand[43]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input107 (.I(b_operand[44]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input108 (.I(b_operand[45]),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input109 (.I(b_operand[46]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input110 (.I(b_operand[47]),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input111 (.I(b_operand[48]),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input112 (.I(b_operand[49]),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input113 (.I(b_operand[4]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input114 (.I(b_operand[50]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input115 (.I(b_operand[51]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input116 (.I(b_operand[52]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input117 (.I(b_operand[53]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input118 (.I(b_operand[54]),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input119 (.I(b_operand[55]),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input120 (.I(b_operand[56]),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input121 (.I(b_operand[57]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input122 (.I(b_operand[58]),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input123 (.I(b_operand[59]),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input124 (.I(b_operand[5]),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input125 (.I(b_operand[60]),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input126 (.I(b_operand[61]),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input127 (.I(b_operand[62]),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input128 (.I(b_operand[63]),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input129 (.I(b_operand[6]),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input130 (.I(b_operand[7]),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input131 (.I(b_operand[8]),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input132 (.I(b_operand[9]),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output133 (.I(net133),
    .Z(ALU_Output[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output134 (.I(net134),
    .Z(ALU_Output[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output135 (.I(net135),
    .Z(ALU_Output[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output136 (.I(net136),
    .Z(ALU_Output[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output137 (.I(net137),
    .Z(ALU_Output[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output138 (.I(net138),
    .Z(ALU_Output[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output139 (.I(net139),
    .Z(ALU_Output[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output140 (.I(net140),
    .Z(ALU_Output[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output141 (.I(net141),
    .Z(ALU_Output[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output142 (.I(net142),
    .Z(ALU_Output[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output143 (.I(net143),
    .Z(ALU_Output[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output144 (.I(net144),
    .Z(ALU_Output[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output145 (.I(net145),
    .Z(ALU_Output[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output146 (.I(net146),
    .Z(ALU_Output[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output147 (.I(net147),
    .Z(ALU_Output[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output148 (.I(net148),
    .Z(ALU_Output[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output149 (.I(net149),
    .Z(ALU_Output[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output150 (.I(net150),
    .Z(ALU_Output[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output151 (.I(net151),
    .Z(ALU_Output[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output152 (.I(net152),
    .Z(ALU_Output[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output153 (.I(net153),
    .Z(ALU_Output[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output154 (.I(net154),
    .Z(ALU_Output[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output155 (.I(net155),
    .Z(ALU_Output[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output156 (.I(net156),
    .Z(ALU_Output[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output157 (.I(net157),
    .Z(ALU_Output[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output158 (.I(net158),
    .Z(ALU_Output[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output159 (.I(net159),
    .Z(ALU_Output[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output160 (.I(net160),
    .Z(ALU_Output[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output161 (.I(net161),
    .Z(ALU_Output[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output162 (.I(net162),
    .Z(ALU_Output[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output163 (.I(net163),
    .Z(ALU_Output[37]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output164 (.I(net164),
    .Z(ALU_Output[38]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output165 (.I(net165),
    .Z(ALU_Output[39]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output166 (.I(net166),
    .Z(ALU_Output[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output167 (.I(net167),
    .Z(ALU_Output[40]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output168 (.I(net168),
    .Z(ALU_Output[41]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output169 (.I(net169),
    .Z(ALU_Output[42]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output170 (.I(net170),
    .Z(ALU_Output[43]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output171 (.I(net171),
    .Z(ALU_Output[44]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output172 (.I(net172),
    .Z(ALU_Output[45]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output173 (.I(net173),
    .Z(ALU_Output[46]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output174 (.I(net174),
    .Z(ALU_Output[47]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output175 (.I(net175),
    .Z(ALU_Output[48]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output176 (.I(net176),
    .Z(ALU_Output[49]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output177 (.I(net177),
    .Z(ALU_Output[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output178 (.I(net178),
    .Z(ALU_Output[50]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output179 (.I(net179),
    .Z(ALU_Output[51]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output180 (.I(net180),
    .Z(ALU_Output[52]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output181 (.I(net181),
    .Z(ALU_Output[53]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output182 (.I(net182),
    .Z(ALU_Output[54]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output183 (.I(net183),
    .Z(ALU_Output[55]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output184 (.I(net184),
    .Z(ALU_Output[56]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output185 (.I(net185),
    .Z(ALU_Output[57]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output186 (.I(net186),
    .Z(ALU_Output[58]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output187 (.I(net187),
    .Z(ALU_Output[59]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output188 (.I(net188),
    .Z(ALU_Output[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output189 (.I(net189),
    .Z(ALU_Output[60]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output190 (.I(net190),
    .Z(ALU_Output[61]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output191 (.I(net191),
    .Z(ALU_Output[62]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output192 (.I(net192),
    .Z(ALU_Output[63]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output193 (.I(net193),
    .Z(ALU_Output[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output194 (.I(net194),
    .Z(ALU_Output[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output195 (.I(net195),
    .Z(ALU_Output[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output196 (.I(net196),
    .Z(ALU_Output[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output197 (.I(net197),
    .Z(Exception[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output198 (.I(net198),
    .Z(Exception[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output199 (.I(net199),
    .Z(Exception[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output200 (.I(net200),
    .Z(Exception[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output201 (.I(net201),
    .Z(Overflow[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output202 (.I(net202),
    .Z(Overflow[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output203 (.I(net203),
    .Z(Overflow[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output204 (.I(net204),
    .Z(Overflow[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output205 (.I(net205),
    .Z(Underflow[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output206 (.I(net206),
    .Z(Underflow[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output207 (.I(net207),
    .Z(Underflow[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output208 (.I(net208),
    .Z(Underflow[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(Operation[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(Operation[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(Operation[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(Operation[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A1 (.I(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__A1 (.I(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__A1 (.I(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__A2 (.I(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__A3 (.I(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A2 (.I(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A2 (.I(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A2 (.I(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__A1 (.I(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__A1 (.I(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A2 (.I(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A1 (.I(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__I (.I(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A2 (.I(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__B (.I(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__B (.I(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A1 (.I(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__A1 (.I(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__B2 (.I(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__A1 (.I(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A1 (.I(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A1 (.I(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__A2 (.I(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A2 (.I(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A2 (.I(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__A2 (.I(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__B2 (.I(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__B (.I(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A3 (.I(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A1 (.I(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A2 (.I(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A1 (.I(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A1 (.I(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06567__A1 (.I(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A1 (.I(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A1 (.I(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A2 (.I(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A2 (.I(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A2 (.I(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A3 (.I(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A1 (.I(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__A1 (.I(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A1 (.I(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__A1 (.I(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A1 (.I(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A2 (.I(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__A1 (.I(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A2 (.I(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__A2 (.I(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A2 (.I(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A1 (.I(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A1 (.I(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__A1 (.I(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A2 (.I(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A3 (.I(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A2 (.I(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A2 (.I(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__A2 (.I(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A2 (.I(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A3 (.I(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__B1 (.I(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__B1 (.I(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__B1 (.I(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A2 (.I(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A2 (.I(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__C2 (.I(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__A1 (.I(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__A1 (.I(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A1 (.I(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A2 (.I(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A2 (.I(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A2 (.I(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A2 (.I(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__B1 (.I(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__B1 (.I(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A2 (.I(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__B1 (.I(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__B1 (.I(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__B1 (.I(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__B1 (.I(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__B1 (.I(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__C (.I(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__A1 (.I(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A1 (.I(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__A1 (.I(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__I (.I(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A1 (.I(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A1 (.I(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A1 (.I(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A1 (.I(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__A1 (.I(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A1 (.I(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A1 (.I(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__A1 (.I(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A1 (.I(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A1 (.I(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__A1 (.I(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__A1 (.I(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__A2 (.I(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A1 (.I(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A1 (.I(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__A1 (.I(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__A2 (.I(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A1 (.I(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A1 (.I(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__A2 (.I(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A2 (.I(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A2 (.I(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__A3 (.I(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__A2 (.I(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__B2 (.I(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A1 (.I(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A1 (.I(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A1 (.I(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A2 (.I(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__A2 (.I(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A2 (.I(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A2 (.I(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__C1 (.I(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__B1 (.I(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__B1 (.I(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__B1 (.I(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A1 (.I(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__A1 (.I(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__A1 (.I(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A2 (.I(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A2 (.I(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A2 (.I(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A2 (.I(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__B2 (.I(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__A1 (.I(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A1 (.I(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A1 (.I(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A2 (.I(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__A2 (.I(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A2 (.I(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__I (.I(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__A2 (.I(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A2 (.I(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A2 (.I(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A2 (.I(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__B1 (.I(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A2 (.I(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__I (.I(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__B1 (.I(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__C1 (.I(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A2 (.I(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A2 (.I(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__C1 (.I(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A2 (.I(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__B2 (.I(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__B2 (.I(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A2 (.I(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__B2 (.I(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__B2 (.I(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__B (.I(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__B2 (.I(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A2 (.I(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A2 (.I(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__I (.I(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A2 (.I(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A1 (.I(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A1 (.I(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__I (.I(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A1 (.I(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__A1 (.I(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__A1 (.I(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A1 (.I(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__A1 (.I(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__A2 (.I(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A1 (.I(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A1 (.I(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A1 (.I(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A2 (.I(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A2 (.I(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A2 (.I(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A1 (.I(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__A1 (.I(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A1 (.I(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A1 (.I(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A2 (.I(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__A1 (.I(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A1 (.I(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A1 (.I(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A1 (.I(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__A1 (.I(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A1 (.I(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A1 (.I(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__A1 (.I(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__A1 (.I(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__A1 (.I(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A1 (.I(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__A2 (.I(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A2 (.I(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__A1 (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__A1 (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A2 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A3 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__A2 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__A1 (.I(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A1 (.I(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__B (.I(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__B1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A1 (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A1 (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A1 (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__A1 (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__C (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__C (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__C (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__C (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__B1 (.I(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A2 (.I(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__B1 (.I(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A2 (.I(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__A1 (.I(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A1 (.I(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__A1 (.I(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A1 (.I(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A2 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A2 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A2 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A1 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A1 (.I(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A1 (.I(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A1 (.I(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__A1 (.I(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__A1 (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__A1 (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A2 (.I(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__A2 (.I(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A1 (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06942__A1 (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__A1 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__A1 (.I(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__A1 (.I(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A2 (.I(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A2 (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__A2 (.I(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A2 (.I(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06942__A3 (.I(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A1 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A1 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__A2 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__A2 (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A2 (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__A2 (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__A2 (.I(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A2 (.I(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A1 (.I(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__A2 (.I(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A1 (.I(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A2 (.I(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07084__A2 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__A2 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__I (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__B2 (.I(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A2 (.I(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A2 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A2 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A1 (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A1 (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A1 (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__A1 (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07073__A2 (.I(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__A2 (.I(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A3 (.I(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__A2 (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__B1 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__B1 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A2 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__I (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A2 (.I(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A2 (.I(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A2 (.I(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A2 (.I(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__C (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__C (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__C (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__C (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__B (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A2 (.I(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__A2 (.I(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A2 (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__A1 (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A2 (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A2 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A2 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A2 (.I(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A2 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A2 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__I (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__A1 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A2 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__A2 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A2 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A3 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__A1 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A1 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A1 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__A1 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__B (.I(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__B (.I(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__B (.I(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__B (.I(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A1 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A1 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A1 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__A2 (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A3 (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__A3 (.I(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__A2 (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A2 (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A2 (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A2 (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A2 (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__I (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__B (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__B (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__B (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__B (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A1 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A1 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A1 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__I (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__B2 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__B2 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A1 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__C1 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__A1 (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A2 (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__I (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A2 (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A1 (.I(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__A2 (.I(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__B (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__B1 (.I(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A4 (.I(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A2 (.I(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__I (.I(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A2 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A2 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A1 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__I (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__B2 (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A1 (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A2 (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A1 (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__I (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A1 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A1 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__A2 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__I (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A1 (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A1 (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A1 (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__I (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A2 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__B2 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A1 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A1 (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A1 (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A1 (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A1 (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A2 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__A2 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A2 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__I (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A2 (.I(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A2 (.I(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__I (.I(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A2 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A2 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A4 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A1 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__B2 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A2 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__I (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__A2 (.I(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__I (.I(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__I (.I(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A1 (.I(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A1 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A1 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__I (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A2 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A1 (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__B2 (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A2 (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__I (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A1 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A2 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__I (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__I (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A1 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A1 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A1 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__I (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A2 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A1 (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A1 (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A1 (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__I (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A2 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__I (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A2 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A1 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__I (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__I (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A1 (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A2 (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__A2 (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__I (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A1 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A2 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A2 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__A1 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A1 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A1 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__I (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A1 (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A1 (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A1 (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__I (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A1 (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A1 (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__I (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__I (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__B2 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A1 (.I(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A1 (.I(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A1 (.I(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__I (.I(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A1 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__A2 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A2 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__I (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A1 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A2 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__A2 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A2 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A2 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__I (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A2 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A1 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__A2 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__I (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A2 (.I(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__A1 (.I(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A2 (.I(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A2 (.I(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A2 (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A2 (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A1 (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__I (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A1 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A1 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A1 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__I (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A2 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A2 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A1 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__I (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A2 (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__I (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A1 (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A1 (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A2 (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A1 (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__A2 (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__I (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A2 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A2 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A1 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__I (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A2 (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__A1 (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A2 (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__I (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A2 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A1 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__A1 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__I (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A2 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A2 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A1 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__I (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A2 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A1 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__I (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__A1 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A2 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A1 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__B1 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__I (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__A2 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A1 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A2 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__I (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A2 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A2 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__B2 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__I (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A1 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__A1 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A1 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A2 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A2 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A2 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__I (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A2 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A2 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A2 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__I (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A2 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A2 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__A1 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__I (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__B2 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A2 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A2 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A2 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__I (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A2 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A2 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A1 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__I (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A2 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A2 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A1 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__I (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__B (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A2 (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__A1 (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__A1 (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A1 (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__I (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A1 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A1 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__A2 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__A2 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A2 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A2 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A2 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__I (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A2 (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__B1 (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A2 (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__I (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A2 (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A1 (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__I (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A2 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__I (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__B1 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A1 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A2 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__I (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A2 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A1 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__A1 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A1 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A2 (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__B (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__I (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__A1 (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__A1 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A1 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A1 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A1 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A2 (.I(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A1 (.I(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__B1 (.I(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__A2 (.I(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A2 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A2 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A1 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__I (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A1 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A2 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__A1 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__I (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__A2 (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A2 (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__I (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__I (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A2 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A2 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__A2 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__I (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A2 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__A2 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__A2 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__B1 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A1 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A2 (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A1 (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__I (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__A2 (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__B2 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A2 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A2 (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A2 (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__I (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A2 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__B2 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A1 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__I (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A2 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A2 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A2 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__I (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A1 (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A1 (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__I (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A1 (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A2 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A2 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__I (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A2 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__B2 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__A2 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__I (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A2 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A2 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__I (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A2 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__C1 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A1 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__A1 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A2 (.I(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A2 (.I(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__I (.I(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__B2 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A1 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A1 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__A1 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A1 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A1 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A2 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A1 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__B2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__A2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__A1 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A1 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A2 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__A2 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A2 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__A2 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A1 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__A2 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A1 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__A1 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A1 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__I (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A2 (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A2 (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__I (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A1 (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A1 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A1 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__I (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A1 (.I(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A1 (.I(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A1 (.I(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__A1 (.I(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__I (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07392__I (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A1 (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__I (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A2 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A2 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A2 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__A2 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__B1 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A1 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A1 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A1 (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A1 (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__I (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A1 (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A1 (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__I (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A1 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A1 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A2 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A2 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A1 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A2 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A2 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A1 (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A2 (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__A2 (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__I (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__A1 (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A1 (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A2 (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__I (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A1 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A2 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__A2 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__I (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__A2 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__A2 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A1 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A2 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A2 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A2 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A2 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__B (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A2 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A2 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A2 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A2 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A2 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__I (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A1 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A1 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A1 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__I (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__A2 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A1 (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A1 (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A1 (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__B2 (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A2 (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__B (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A1 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A3 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__B2 (.I(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__B1 (.I(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__B1 (.I(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A2 (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A3 (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A1 (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__B1 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A2 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A1 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A1 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A1 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__B (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A2 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A2 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A2 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A2 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__B2 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A1 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A1 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A1 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__B1 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__B1 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__C1 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__B1 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__S (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A1 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__S (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A2 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A1 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A1 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A1 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A1 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A2 (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A2 (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A2 (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__B1 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__B1 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A2 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__B1 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A2 (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__A2 (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__B1 (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A2 (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__B2 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A3 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__B2 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__B2 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A1 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A1 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A1 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__A1 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A1 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A1 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A4 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__I (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A3 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A3 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A1 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A1 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__B2 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__B2 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__B2 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__B2 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A2 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A2 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__A2 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__I (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A2 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A2 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A2 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A1 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__B1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A2 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__B2 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__B2 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__B2 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__B2 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__C (.I(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A2 (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__A2 (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__B (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__I (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A2 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A2 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__I (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__A1 (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__A1 (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A1 (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A1 (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A2 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A3 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__I (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A2 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A1 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A1 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A1 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__B2 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A1 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A1 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__A1 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A2 (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A2 (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__A1 (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__I (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A2 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A2 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A2 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__B1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__A2 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A2 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__B1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A2 (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A2 (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__I (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__A1 (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A1 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A1 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__A1 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__C1 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__I (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05677__I (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A2 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A2 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A3 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A1 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__I (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A2 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A2 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A2 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A2 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__A1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__B1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A3 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A2 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A2 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A2 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__A1 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A1 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__I (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05678__I (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A2 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__A1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A2 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__A2 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A2 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__B1 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__A2 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05679__I (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A1 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A1 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__A1 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__B1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A3 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__B (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__B2 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__B2 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__B2 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A2 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A2 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A3 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A2 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05697__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05692__I (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05681__I (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A1 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A1 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__B (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__S (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__B (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__B (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__B (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__B (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A2 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__A2 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__A2 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__A2 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A2 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A2 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A1 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__I (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A2 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A2 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A2 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__A1 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A3 (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__A2 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A2 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A2 (.I(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A2 (.I(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__A3 (.I(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__A2 (.I(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__B2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__A1 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__I (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A1 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__B1 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__B1 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__B1 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__B1 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__A1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__B1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A3 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A3 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__C2 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__B2 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A1 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A1 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A1 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A1 (.I(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A1 (.I(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A1 (.I(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__B1 (.I(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A1 (.I(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A2 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05690__I (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__B2 (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__A2 (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A1 (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__A3 (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A1 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A1 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A1 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__A2 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A2 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05691__I (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A1 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A1 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A2 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A2 (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A2 (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__I (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05754__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__B (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__A2 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A2 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A2 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__A2 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__B2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__B2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__B2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__B2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A1 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A1 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A1 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__A2 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A2 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A2 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__B1 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__B2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__I (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__B1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__B2 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__C2 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__C2 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__B2 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__A2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__B2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__A2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__A1 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__B1 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A1 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__B (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__I (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__B2 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A3 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A1 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A1 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A1 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__A2 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05737__I (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05695__A2 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__A1 (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__A2 (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A1 (.I(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A2 (.I(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A1 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__A1 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A1 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__A1 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A1 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A2 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__A1 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A1 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A1 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A1 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05697__A2 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A1 (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A1 (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A1 (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A2 (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A3 (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__A3 (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__B (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A1 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A1 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A1 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__I (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A1 (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A1 (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A1 (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__I (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A1 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A1 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A2 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__I (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__B2 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__A1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A2 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A2 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A2 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__C1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A1 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A1 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A1 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A1 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__I (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05742__I (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05701__A2 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__B2 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__B (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A3 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__A1 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__B1 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__B1 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__B1 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05703__I (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A1 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A1 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A2 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A3 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__A1 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__B1 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__B1 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05714__A1 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A2 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A2 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__B1 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A1 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__B2 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A2 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A3 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A1 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__A1 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A3 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__B (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__B1 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__B2 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__B2 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__B2 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__B2 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__B1 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A1 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__A2 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A3 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__A2 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A1 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A1 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A1 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A1 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A2 (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A2 (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A2 (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A2 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A2 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__B1 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__B1 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__I (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__I (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05714__A2 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A1 (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A3 (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A2 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A2 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A1 (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A1 (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A2 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__A2 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A2 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A3 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__A1 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05741__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05712__A4 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__I (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__I (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__I (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05713__I (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A2 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__B2 (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__B (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A1 (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__B (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__I (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__I (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05714__A3 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A2 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__I (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__I (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__C1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__B1 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A1 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__B (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05715__B (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__B2 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A2 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A2 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A2 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__B2 (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__B (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A3 (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A1 (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__B1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__A2 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__B2 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__I (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__B2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__B2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__A2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05719__I (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A2 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A2 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A2 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A3 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__B (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A1 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__A1 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A1 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__I (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A2 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A2 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A3 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A2 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A3 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__B1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__B2 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__B2 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__C2 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A3 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A2 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A2 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A1 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05723__I (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__B (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__I (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A1 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__A1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A2 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A2 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A1 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A1 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A2 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A2 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A2 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A3 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__A2 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__A2 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05729__I (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A2 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__B2 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__A2 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__I (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05731__A2 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__B1 (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A3 (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__B (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__A1 (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__B2 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A1 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A1 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A1 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A1 (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A1 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__I (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__I (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__I (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__A2 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A1 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A1 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A2 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__I (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__I (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__I (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__I (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A1 (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A2 (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A3 (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A2 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__B1 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__B1 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__B1 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__A1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A2 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05954__I (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05738__I (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A2 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A2 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A2 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__B (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__I (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A1 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__A2 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__B2 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05751__A1 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A1 (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A1 (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A2 (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__A1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__A1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__A1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A1 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A1 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__I (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__I (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__C2 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__A2 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A1 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A2 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A1 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A2 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A1 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A1 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A1 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A2 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A2 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A1 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A1 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__A2 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__A2 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A2 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A2 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__A3 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__A3 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A2 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A2 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A2 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A2 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A2 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__B1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__C (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05750__A2 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__C2 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A2 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A2 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05751__A2 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A2 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A2 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A1 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A2 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A2 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A2 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A3 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A1 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A1 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__I (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__I (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__A2 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A2 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A2 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__C (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__A2 (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A2 (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A3 (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__A3 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A3 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__B (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A2 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__C (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__B (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__B (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A1 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A2 (.I(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A2 (.I(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A1 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A1 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A2 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__A2 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__A2 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__A2 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__I (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A1 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A1 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A2 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A2 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A2 (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__A2 (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__A2 (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__I (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A2 (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A2 (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A2 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A4 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__A2 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A2 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A2 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A1 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A2 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A2 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A2 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A1 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A1 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A2 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A2 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A2 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__A2 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A2 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A2 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A3 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A1 (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__C (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A1 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__B2 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06915__A2 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05766__I (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A2 (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__B1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__I (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A1 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__I (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__A1 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A2 (.I(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__I (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__I (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A2 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__A2 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__A2 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A1 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__A2 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A2 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A2 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A2 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A2 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__A2 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A2 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A2 (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A1 (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__I (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__I (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__A1 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A2 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__B2 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__A1 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__A1 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A2 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A2 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A3 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A2 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A1 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A2 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A2 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__A2 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__I (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__A2 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__B (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A2 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A3 (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__A1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__I (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__A2 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A1 (.I(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A1 (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A1 (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__A2 (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A3 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A2 (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__I (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A1 (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__I (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A2 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A3 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A3 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__A3 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A3 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A2 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A2 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A1 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A1 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A1 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A1 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__I (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__I (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A1 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A1 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A1 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__I (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__I (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A1 (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A1 (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A1 (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__C1 (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__I (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A2 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__I (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A2 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A2 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A2 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__A2 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__I (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A2 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__I (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A2 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__I (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__B2 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A2 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__I (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05783__I (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__C2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__B1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A2 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A2 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A2 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__I (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__B2 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A2 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__B2 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A1 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A1 (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A1 (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__I (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A4 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__I (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__I (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__B2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__B2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__A2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__I (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__B1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__B1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__A2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__B2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__I (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__A1 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A1 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__I (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A2 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__B (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A2 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__I (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__I (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A1 (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A1 (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__I (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__A1 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A2 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A2 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__I (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05786__I (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__I (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__I (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A2 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__I (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A1 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A1 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A1 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__A1 (.I(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__B2 (.I(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A2 (.I(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A2 (.I(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A1 (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__I (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A1 (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A1 (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__A1 (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A1 (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__A2 (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__I (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__I (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__I (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__I (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__B2 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A2 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A2 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__I (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__I (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A1 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A1 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__I (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__I (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__A1 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A2 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A1 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__B1 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A2 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__I (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06675__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A2 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__I (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__I (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__A1 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__A1 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A2 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__I (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A1 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A1 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__I (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A1 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A1 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A1 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__I (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__I (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A1 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A1 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A1 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__I (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A1 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__B1 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__I (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A2 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__A2 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__B2 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A2 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__B2 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A2 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__A2 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A2 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A1 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__I (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A2 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A2 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A2 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__A2 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A2 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__B1 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A2 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__I (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__I (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A1 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A1 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__I (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A2 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__B1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A2 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__A2 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A1 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A2 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__I (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A1 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__I (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05923__A2 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__I (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A2 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__I (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A1 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__I (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A2 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__I (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A2 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__I (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__A2 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A3 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__I (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__I (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A2 (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A1 (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A1 (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__I (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A1 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__I (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A2 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A3 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__I (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__I (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__B1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A2 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__I (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A2 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A1 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__I (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__A2 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A3 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A1 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A1 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__I (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A2 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__I (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__I (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A2 (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A3 (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__I (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__I (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A2 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A1 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__I (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A2 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A2 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A2 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A1 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__I (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__B1 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A4 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__I (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A2 (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A2 (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A1 (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__I (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A1 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__I (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__I (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A2 (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A1 (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__I (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__I (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A2 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A3 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A2 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__I (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A1 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A2 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__I (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A2 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__B1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__B1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A2 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A1 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A1 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__I (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A2 (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A2 (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A1 (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__I (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__I (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A2 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A1 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__B1 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__I (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__A2 (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A2 (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A1 (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__I (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A2 (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A2 (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A1 (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__I (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A2 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__I (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A1 (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__A2 (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__I (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05796__I (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__B2 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__I (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A2 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__B2 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__B2 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__B2 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A2 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A2 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A2 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A2 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__I (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__I (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__I0 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A2 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__I (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__I (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A2 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09344__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__I (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__I (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__B (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__B1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A2 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A2 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__B2 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A2 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__I (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__B (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A2 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A3 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A1 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A1 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__A2 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__B2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A1 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A1 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A1 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__B1 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A1 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__A2 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__A2 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05800__I (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A1 (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__I (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__I (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A2 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A1 (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A3 (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A2 (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__I (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__A1 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__B1 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__I (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A1 (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A2 (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__B (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__I (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__I (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A2 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A2 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__I (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A2 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__I (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__I (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A2 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A1 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__B2 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A3 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A1 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__B2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__B2 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__I (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A4 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A1 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A1 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A1 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A1 (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A1 (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A1 (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A1 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A2 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__I (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A2 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__I (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A2 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__B (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__I (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A3 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__I (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A2 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__B (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__I (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A4 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__B (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__I (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__C (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A2 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05808__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A1 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__I (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__I (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__I (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A2 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__A4 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__I (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A1 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__I (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__I (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A1 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__B1 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A1 (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A2 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__B1 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A2 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A2 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__B2 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A2 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A2 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A2 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__I (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A2 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__I (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A1 (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A2 (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A2 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A2 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__B2 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__B1 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__I (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__A2 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A2 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A2 (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A2 (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__I (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__I (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A2 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A2 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__I (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A2 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A3 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__I (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__I (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__B1 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A2 (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A3 (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A2 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__A2 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__A1 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A1 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__I (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A2 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A2 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A2 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__I (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__A2 (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A2 (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A1 (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A1 (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__B2 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A2 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__A2 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__A1 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A1 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__I (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A2 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A2 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A2 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__B2 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__B2 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__C2 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__B1 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__B1 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A1 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__B2 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A2 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A2 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__I (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A2 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A2 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A3 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A3 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A3 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A3 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A4 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A3 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__A2 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__I (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A2 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__B1 (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__B2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__B2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__B2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__B2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__A2 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__B1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__I (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A1 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A1 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A1 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A1 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__A2 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A2 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A1 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05816__I (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__B (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A4 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A2 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A1 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A2 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__I (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A2 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__B2 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__I (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__A2 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A2 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A2 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A2 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__B2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A2 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A1 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A1 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__C1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__I (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A2 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__S (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A3 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__A2 (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__A1 (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__A1 (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__I (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A2 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A2 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A1 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__B1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A2 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A2 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A2 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A4 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A2 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__A1 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__A2 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A3 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A4 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A4 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A4 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A2 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__I (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__I (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A3 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__B2 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A3 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A2 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__B1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__B2 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__B2 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__B1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A2 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__B2 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A2 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__S (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__S (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A3 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__I (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A2 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A2 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A2 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A2 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A2 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A2 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__A2 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A1 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A1 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A4 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A2 (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A2 (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__B1 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A2 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A2 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A2 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A2 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A3 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__A2 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A2 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A2 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__I (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__B2 (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__B2 (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__B2 (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A2 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A3 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__B1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A2 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A2 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__A2 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__I (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__A2 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A2 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__I (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A3 (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A1 (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A1 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A1 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A2 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__I (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A1 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A1 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A1 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A1 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__A1 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__B (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__C2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__A1 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__A1 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__A1 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A1 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A1 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A1 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A1 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A1 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__B2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A4 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A4 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A4 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A1 (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__I (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A2 (.I(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__A1 (.I(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A3 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__A3 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A2 (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A2 (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A2 (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__I (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A2 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A3 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A1 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__B1 (.I(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__B2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__B2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__B2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A2 (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A1 (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A1 (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__A3 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__B2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05837__I (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__C (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__B (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__B (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__A1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__A1 (.I(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__A1 (.I(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A1 (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A1 (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A2 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__A2 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__A1 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__I (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A4 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__B2 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A2 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__A3 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A2 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A2 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A2 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__I (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__I (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__C1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__I (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__A2 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__A3 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A2 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__B1 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A1 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__I (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A1 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A1 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A2 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__A1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__I (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A3 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__A1 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A1 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A1 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A2 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A2 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A2 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A1 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A3 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A3 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A2 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A2 (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A2 (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A4 (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A2 (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A2 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__A2 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A2 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__I (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__A4 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__I (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__I (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__A2 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A3 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__I (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A2 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__B1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__I (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__I (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A2 (.I(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A2 (.I(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__A2 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__A2 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A2 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05853__A2 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A2 (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A1 (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__B2 (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__B2 (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__B1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A1 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__A2 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A2 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A2 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A1 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A2 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A1 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__A1 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A1 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__B (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__A2 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A1 (.I(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A1 (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A1 (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A2 (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__B2 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A1 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__I (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A2 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__A2 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__I (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__A2 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__B (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A1 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A1 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__B2 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A1 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__B2 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A1 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A2 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A1 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__B2 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__B (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A1 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A1 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06100__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A1 (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__B1 (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__A2 (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A1 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A1 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__B2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A2 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A2 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A2 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A1 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A3 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__A1 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A2 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A4 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A1 (.I(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__B1 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__A1 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A2 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A2 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A2 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A1 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A1 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A1 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A3 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A2 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A1 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__B (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A3 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A1 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A1 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A2 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A2 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A3 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__A2 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A2 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__I (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__B1 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__A2 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__A2 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__I (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__B (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A1 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A2 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A2 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__A2 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A1 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__A1 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__I (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A3 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A2 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A2 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__I (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__I (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__B2 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A1 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A2 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A2 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__B (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__B1 (.I(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__A1 (.I(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A2 (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A2 (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__B (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__B (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A1 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__B (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A2 (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A2 (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__A1 (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__I (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A3 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A2 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A2 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A1 (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A1 (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A2 (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__A1 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__B2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A1 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A1 (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A2 (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A1 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A3 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__B1 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A2 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__B (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A2 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__B (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__I (.I(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__B2 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__A1 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__A1 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__A1 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A1 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A1 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A1 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A2 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A2 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A1 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A1 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A3 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A2 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A2 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A2 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A2 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A2 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A2 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A3 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A2 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__C2 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A2 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A1 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__I (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__I (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__A1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A2 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__B2 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A1 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__I (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A2 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A2 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__B2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__I (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A1 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__A1 (.I(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A1 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__A1 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A2 (.I(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A2 (.I(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A2 (.I(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A3 (.I(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A1 (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A1 (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__A2 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A1 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A1 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__I (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A2 (.I(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__B1 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A2 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__B2 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A2 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__I (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A1 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A2 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A1 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A1 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A4 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A2 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A2 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__B2 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__I (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A2 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__I (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A2 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__I (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A1 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A2 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A2 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__B1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__A1 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A1 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A3 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__A2 (.I(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A2 (.I(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A3 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__B (.I(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A2 (.I(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A1 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A1 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__I (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A1 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A2 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A1 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A1 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__B (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A1 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A1 (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__I (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A2 (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__I (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A1 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A1 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__A2 (.I(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A2 (.I(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__B2 (.I(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__A1 (.I(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__A1 (.I(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__I (.I(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__B (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__A1 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A1 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A2 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__A3 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A1 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A1 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A1 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A2 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A2 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A2 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A2 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__I (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A2 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A2 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__I (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__B (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__I (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A1 (.I(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A2 (.I(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A2 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__A2 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A2 (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A2 (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A1 (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A1 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A1 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A2 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A1 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__A1 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A1 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__A1 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__A1 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A1 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A1 (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A1 (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A2 (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__I (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__A2 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__A1 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09924__A1 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__A2 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09924__A2 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__B (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A1 (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A2 (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__A2 (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__A2 (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A1 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A1 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__A1 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__I (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A1 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__A2 (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A3 (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A1 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A1 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A1 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__I (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A2 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__I (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__A1 (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A2 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A2 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A3 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__B (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__C (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A1 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A2 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A2 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A2 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__B (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__A2 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A2 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__A1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__A3 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A3 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A3 (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__I (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__I (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__B1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__B2 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__B2 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__I (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__B1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A4 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A2 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__I (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__I (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__C2 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__B1 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A2 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A1 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__I (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__I (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__I (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__B2 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__I (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__I (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A1 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A1 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A1 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__I (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__A1 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A2 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A2 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__I (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__I (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__B2 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A2 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A1 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__C2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A1 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A1 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__A2 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A2 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__I (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__I (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A2 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__A2 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A2 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__I (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__A2 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A2 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A2 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__I (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A2 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A2 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A2 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A2 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A2 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__A2 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__I (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__I (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A1 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__I (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__I (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A1 (.I(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__A1 (.I(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A1 (.I(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__I (.I(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A1 (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A1 (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A2 (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__I (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A2 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__I (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A2 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__I (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__I (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__A1 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A2 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A2 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__B1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__I (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A1 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__I (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A1 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A1 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__I (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A1 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A2 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__I (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__I (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__A1 (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A2 (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A2 (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A1 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A1 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__I (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__A1 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A1 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__A2 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__I (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__B2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__I (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__I (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A1 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A1 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__A1 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__I (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__I (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__I (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A1 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__B1 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A1 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__I (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A1 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__I (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__A2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__A2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A2 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A1 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__A1 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__I (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__I (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A2 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A2 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A2 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__I (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__A2 (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__I (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A2 (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A2 (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A2 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__I (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__A2 (.I(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A2 (.I(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A2 (.I(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__I (.I(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A2 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A2 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__I (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A1 (.I(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A1 (.I(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A1 (.I(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A1 (.I(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__B2 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A1 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__A1 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__I (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A1 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A1 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A2 (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__A2 (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__I (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__I (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__B2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__I (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__I (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__B2 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__I (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A2 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__B2 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__I (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__A1 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__I (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__A1 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__A1 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__I (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__B2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__I (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__I (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__A2 (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__A2 (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A1 (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__I (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__B1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__I (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A2 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__I (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A2 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A2 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A2 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A1 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__I (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__B1 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A1 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__A1 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__I (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A2 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__A2 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__I (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A1 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__B2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__A2 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__I (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__A2 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__I (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A2 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__I (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__I (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A2 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A3 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A2 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__I (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__A2 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__I (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A1 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__I (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A1 (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A1 (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A2 (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__I (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__I (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__B (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A2 (.I(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__I (.I(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__A1 (.I(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__I (.I(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__A2 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A2 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__I (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A2 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A2 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A1 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__I (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__I (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A2 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__A2 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A2 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__I (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__I (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__B1 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__A2 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__A2 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__I (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__I (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A2 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A2 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__I (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A2 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A1 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A1 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A1 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A2 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__B2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__B2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__B2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A2 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A2 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A2 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__I (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__A2 (.I(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A2 (.I(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__I (.I(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__I (.I(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__A4 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__I (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__B1 (.I(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A1 (.I(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__A1 (.I(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__I (.I(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__A2 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A2 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A2 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__I (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__I (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__I (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__B1 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__B (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__B (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__I (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__A2 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A2 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__A1 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A1 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A1 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__B (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__C2 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A1 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A1 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__I (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__A1 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__A1 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A2 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__I (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A1 (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__A1 (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__A1 (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A1 (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A1 (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A1 (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__A1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A1 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A1 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__I (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A2 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__B1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__I (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__I (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__B (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__I (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__A1 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__B2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__I (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A1 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A1 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__A2 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__I (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__A1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__I (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__I (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__A2 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__I (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__I (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__A3 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A1 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__C (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__A2 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__A1 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A1 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A2 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__I (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A1 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A1 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__I (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__I (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A1 (.I(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A1 (.I(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A2 (.I(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__I (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__I (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A1 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__B2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A1 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A1 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__B2 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__A1 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__A1 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A2 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__B (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__I (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A3 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__I (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__B (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__A1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A2 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__B (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__I (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A3 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__I (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__I (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__B (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__B (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__I (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__I (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__B1 (.I(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A2 (.I(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A3 (.I(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A2 (.I(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__A1 (.I(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A1 (.I(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A1 (.I(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A2 (.I(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__I (.I(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A3 (.I(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A3 (.I(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__A2 (.I(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__A2 (.I(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__B2 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A2 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__B (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A3 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__B1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__I (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__I (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__I (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__I (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__B2 (.I(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A2 (.I(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__A1 (.I(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A1 (.I(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A1 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__B2 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__A1 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A2 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A2 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A2 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A1 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A1 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A1 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__A1 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__B2 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A1 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A1 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A1 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A3 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A1 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A1 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A1 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A2 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__A1 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__A3 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A2 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__B1 (.I(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__B1 (.I(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A2 (.I(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__B (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__B1 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A2 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__B (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__B1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A2 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__A1 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__A1 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__A2 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A2 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__A1 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__A1 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__B1 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__I (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__I (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A2 (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__I (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__I (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A2 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A2 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A3 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__A1 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A1 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__A2 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A1 (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A1 (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A1 (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__I (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__I (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__I (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__I (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__I (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A2 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__A1 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__B1 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A2 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__A1 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A1 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__B1 (.I(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__B1 (.I(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__I (.I(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__I (.I(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__B1 (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A2 (.I(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__A2 (.I(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A2 (.I(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__A2 (.I(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__B2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__B1 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__B2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__B2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A1 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__A3 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__B1 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__A2 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__B2 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A2 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A2 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__A1 (.I(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A2 (.I(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__A1 (.I(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A2 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A1 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A1 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__I (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A2 (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A2 (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__B2 (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__I (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__B2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A2 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__A2 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A3 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A1 (.I(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__A2 (.I(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__A2 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A2 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__A3 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A2 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A2 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A2 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__I (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A2 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__C1 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A2 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__I (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__I (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A2 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__A3 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__B2 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A1 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A2 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A1 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A1 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__C1 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__B1 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A2 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__A2 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A2 (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__A2 (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__B (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__B (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__B (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__B (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A2 (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__A2 (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A2 (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__I (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A2 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A2 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__A2 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A2 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__A2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__A1 (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__B1 (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A1 (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__C2 (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__A1 (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__A1 (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A1 (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__A1 (.I(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__A2 (.I(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A2 (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A2 (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A2 (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__A1 (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__A2 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A2 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__A2 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__A2 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__B2 (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__A2 (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A1 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__A3 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__I (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__I (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__I (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__I (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__A1 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10569__A1 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A2 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A2 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A2 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__I (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A2 (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__A2 (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__I (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__B1 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A2 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A2 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__B2 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__A2 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__A3 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__I (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__B1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A1 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__A1 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A1 (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A1 (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A2 (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__A1 (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A1 (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__B (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A1 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A1 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__A1 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__A1 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__C (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__I (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__I (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__I (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A2 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A2 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__B1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A2 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__A2 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__A2 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__B (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__B (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__C (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__I (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__A1 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__A3 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A1 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__B2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__B2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__A1 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__A1 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__A1 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__I (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__A1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__B1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__A2 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__B2 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__B (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__B (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A1 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A1 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__A2 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A1 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A1 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A3 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__B (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__B2 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__A2 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A2 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__B1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__A2 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__B2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A3 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A2 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__A2 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A3 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A1 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__A2 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A2 (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A1 (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__A1 (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__B2 (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A2 (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__B2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A1 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A1 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__I0 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A2 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A3 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__B2 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__A1 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A1 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A1 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__A1 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__B2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A1 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A1 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A1 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__A1 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__A1 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__B (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A1 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A1 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__A1 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A1 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A1 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__A1 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A2 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__A2 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A1 (.I(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__A1 (.I(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A1 (.I(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__A1 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__A1 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A2 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A1 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A3 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__A1 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A1 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__B1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__A2 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__A1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A2 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A2 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A2 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A3 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A2 (.I(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A2 (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__B1 (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__B2 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__B (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A2 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A1 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A2 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__A1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__A1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A1 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__A1 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__B (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__B2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__B (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__I (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__A1 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A1 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__B2 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__B2 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__B2 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__B2 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A1 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__B (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A1 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__A1 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__A1 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__B1 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__I (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A2 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A2 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__B1 (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A1 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A3 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__B1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__A2 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A2 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A2 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__A3 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A2 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A1 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A1 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A1 (.I(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A1 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A1 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__A2 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A3 (.I(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A1 (.I(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A1 (.I(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A1 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A1 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A2 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A1 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__B (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__S (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__I (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A2 (.I(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A2 (.I(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A2 (.I(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A1 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__S (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__S (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A2 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A1 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A1 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A2 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A1 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A3 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A1 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__S (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__B (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__A2 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__A2 (.I(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__A2 (.I(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A2 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A1 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__B (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__B (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__B (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__A1 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__A1 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A2 (.I(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__A1 (.I(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__A1 (.I(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A1 (.I(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__B1 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__A1 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A1 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A1 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__A2 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A3 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__A1 (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__A1 (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A1 (.I(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__A2 (.I(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__B2 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__A2 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A1 (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A1 (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__B2 (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A2 (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__B2 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__B2 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__A2 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__A1 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A1 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A1 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__A1 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__C (.I(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__A1 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A1 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A2 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A2 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A2 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A1 (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__A2 (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A2 (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A1 (.I(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A2 (.I(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A3 (.I(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A1 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__A1 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__A1 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__A1 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__A2 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A1 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__A2 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__A2 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A2 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A2 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__A3 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__A3 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A2 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__A2 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A1 (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A1 (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__I (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06030__I (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__A1 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A1 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A1 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A1 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A1 (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A1 (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A2 (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__A1 (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__B (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__A2 (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A1 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A1 (.I(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A1 (.I(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A2 (.I(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A2 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__A1 (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A2 (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__A1 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A1 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__A2 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A2 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A1 (.I(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A1 (.I(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A2 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A2 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__A2 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A2 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A2 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A1 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A1 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A1 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A2 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A2 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A2 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A2 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A1 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__A2 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__A1 (.I(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__A2 (.I(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A2 (.I(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__I (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A2 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A2 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__I (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__A1 (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__B1 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__A1 (.I(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__A1 (.I(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__I (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__I (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__I (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__I (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11297__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A2 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A2 (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A2 (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A3 (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__A1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__B2 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A2 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__B1 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A2 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A2 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__B (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__A1 (.I(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__A1 (.I(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__B (.I(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A1 (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A1 (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A2 (.I(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A2 (.I(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A1 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__A2 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__A1 (.I(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__A1 (.I(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A2 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A2 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A1 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A2 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A2 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A2 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A2 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__I (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__A1 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__A1 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A3 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__A2 (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__A2 (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__I (.I(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A2 (.I(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__A1 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__A1 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__A2 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A2 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__A2 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A2 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__I (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A1 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__A1 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__A1 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A3 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A2 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A1 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A1 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__B1 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__A2 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__B (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__B (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__B (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__B (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__A1 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A2 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__A1 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A3 (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__B1 (.I(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__B1 (.I(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__B1 (.I(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__C1 (.I(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A3 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A2 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__A2 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__I (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__I (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__I (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__I (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A2 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A2 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A2 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__A2 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__I (.I(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__I (.I(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__I (.I(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__I (.I(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__B2 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__B2 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A3 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__B2 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__B (.I(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__I (.I(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__B (.I(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__I (.I(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A1 (.I(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__B (.I(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__B (.I(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__B (.I(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__B (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A1 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__A1 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__A1 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A1 (.I(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A1 (.I(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__A1 (.I(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__A2 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A2 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__A2 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A2 (.I(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__A2 (.I(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__A3 (.I(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__A2 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__B2 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__B2 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__B2 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__B2 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__C2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__A1 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__A1 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A2 (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__I (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__A2 (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__I (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__B2 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__B2 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A2 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__B2 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__B1 (.I(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__B1 (.I(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__B1 (.I(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__B1 (.I(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A2 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A2 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A1 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__I (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__A2 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A2 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__A2 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A1 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A2 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A2 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A2 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A2 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A2 (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A2 (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__I (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__A1 (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A1 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__A1 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06163__A1 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__B1 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__B2 (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__B2 (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__B2 (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__B2 (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__B1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__C1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__C1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__C1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__C1 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__A3 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__A1 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A1 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__I (.I(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A1 (.I(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__I (.I(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__A1 (.I(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A2 (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A2 (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A2 (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__I (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A2 (.I(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A2 (.I(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A2 (.I(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__A2 (.I(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__B1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__A1 (.I(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__B (.I(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A1 (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__A1 (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__A2 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A2 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__A2 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A1 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__I (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__A1 (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__A1 (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__A2 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A1 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A1 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A1 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A2 (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__A2 (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A3 (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A2 (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__B1 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__I (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__I (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__B1 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__I (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__I (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__I (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__B1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__B (.I(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__A2 (.I(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__I (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A2 (.I(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A2 (.I(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A1 (.I(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I (.I(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__B1 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A2 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A1 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__A1 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__A2 (.I(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__B1 (.I(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A2 (.I(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A1 (.I(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A2 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A2 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A2 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A2 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A1 (.I(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A2 (.I(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__A1 (.I(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__B2 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__A2 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A2 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A2 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__A3 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__A2 (.I(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__B2 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A1 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A1 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A1 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A2 (.I(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__A2 (.I(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A2 (.I(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A2 (.I(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A2 (.I(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__B2 (.I(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__B2 (.I(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__B2 (.I(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__A1 (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__A1 (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A1 (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__B1 (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__I (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__I (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A1 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__I (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__B (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__I (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__I (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__A1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__A1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06344__A1 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A1 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__A1 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A1 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__B1 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A1 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A2 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A2 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A1 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A1 (.I(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A1 (.I(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A2 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A2 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__B1 (.I(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__B2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__B2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__B2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__B2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A2 (.I(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A2 (.I(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A2 (.I(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A2 (.I(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__I (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__I (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__I (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__I (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__B2 (.I(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__B2 (.I(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__B2 (.I(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__B2 (.I(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__B1 (.I(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__B1 (.I(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__A2 (.I(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A2 (.I(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__B1 (.I(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__B1 (.I(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__B1 (.I(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__B1 (.I(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__B2 (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__A1 (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A1 (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A1 (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A2 (.I(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A2 (.I(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A2 (.I(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A2 (.I(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__C2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__C2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__B1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__B1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__B2 (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__A2 (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__A2 (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__I (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__A1 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__B2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A2 (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A2 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A2 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A2 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A2 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__B1 (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__B1 (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__B1 (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__B1 (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A1 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__A1 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A1 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__A1 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__B (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__A3 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A1 (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__S (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__A2 (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A2 (.I(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__A2 (.I(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A1 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A2 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A1 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__A1 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06344__A2 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__A1 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A1 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A1 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__A1 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A2 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__A2 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06427__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A1 (.I(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A1 (.I(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__A2 (.I(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__A2 (.I(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__A1 (.I(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A2 (.I(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__B1 (.I(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A1 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__B2 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__B1 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__B1 (.I(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__B1 (.I(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__B1 (.I(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__B2 (.I(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A2 (.I(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A2 (.I(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__C2 (.I(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__C (.I(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__C2 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A1 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A1 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A1 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A2 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A2 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A2 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A2 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__B1 (.I(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__B1 (.I(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__B1 (.I(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__B1 (.I(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__B1 (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__B1 (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__I (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__B1 (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__C (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A1 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__A2 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A2 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A3 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A1 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A1 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A2 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A2 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A2 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__A1 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A1 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A2 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__I (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__A2 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__B1 (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A2 (.I(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A2 (.I(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A2 (.I(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A2 (.I(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__B2 (.I(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__B2 (.I(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__B2 (.I(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__B2 (.I(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A1 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A1 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__A1 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A1 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A1 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__A2 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A3 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__I (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__B (.I(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__B (.I(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__B (.I(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__B (.I(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A1 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A1 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__A1 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A1 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__A1 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A1 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(a_operand[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(a_operand[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(a_operand[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(a_operand[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(a_operand[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(a_operand[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(a_operand[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(a_operand[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(a_operand[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(a_operand[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(a_operand[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(a_operand[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(a_operand[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(a_operand[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(a_operand[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(a_operand[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(a_operand[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(a_operand[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(a_operand[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(a_operand[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(a_operand[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(a_operand[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(a_operand[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(a_operand[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(a_operand[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(a_operand[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(a_operand[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(a_operand[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(a_operand[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(a_operand[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(a_operand[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(a_operand[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(a_operand[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(a_operand[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(a_operand[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(a_operand[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(a_operand[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(a_operand[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(a_operand[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(a_operand[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(a_operand[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(a_operand[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(a_operand[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(a_operand[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(a_operand[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(a_operand[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(a_operand[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(a_operand[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(a_operand[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(a_operand[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(a_operand[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(a_operand[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(a_operand[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(a_operand[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(a_operand[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(a_operand[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(a_operand[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(a_operand[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(a_operand[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(a_operand[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(a_operand[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(a_operand[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(a_operand[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(a_operand[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(b_operand[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(b_operand[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(b_operand[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(b_operand[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(b_operand[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(b_operand[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(b_operand[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(b_operand[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(b_operand[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(b_operand[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(b_operand[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(b_operand[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(b_operand[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(b_operand[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(b_operand[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(b_operand[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(b_operand[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(b_operand[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(b_operand[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(b_operand[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(b_operand[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(b_operand[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(b_operand[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(b_operand[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(b_operand[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(b_operand[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(b_operand[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(b_operand[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(b_operand[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(b_operand[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(b_operand[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(b_operand[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(b_operand[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(b_operand[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(b_operand[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(b_operand[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(b_operand[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input106_I (.I(b_operand[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input107_I (.I(b_operand[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input108_I (.I(b_operand[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input109_I (.I(b_operand[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input110_I (.I(b_operand[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input111_I (.I(b_operand[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input112_I (.I(b_operand[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input113_I (.I(b_operand[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input114_I (.I(b_operand[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input115_I (.I(b_operand[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input116_I (.I(b_operand[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input117_I (.I(b_operand[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input118_I (.I(b_operand[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input119_I (.I(b_operand[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input120_I (.I(b_operand[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input121_I (.I(b_operand[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input122_I (.I(b_operand[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input123_I (.I(b_operand[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input124_I (.I(b_operand[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input125_I (.I(b_operand[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input126_I (.I(b_operand[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input127_I (.I(b_operand[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input128_I (.I(b_operand[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input129_I (.I(b_operand[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input130_I (.I(b_operand[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input131_I (.I(b_operand[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input132_I (.I(b_operand[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05704__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05684__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05685__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05699__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05683__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05709__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05682__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05676__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05716__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05785__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05776__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__B2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07568__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__B2 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__B2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A2 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A2 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A3 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A3 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A3 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A2 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A2 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A1 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A2 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05696__I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05693__I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A2 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A2 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A2 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__A2 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__A2 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A2 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A2 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A2 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A2 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05906__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05773__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A2 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__A2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A2 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A2 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A2 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A2 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__A1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__A1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A2 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A2 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A2 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A2 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A2 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A2 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A2 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__B2 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__A1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A2 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__A1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A1 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A1 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__A2 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output133_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output134_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output135_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output136_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output137_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output138_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output139_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output140_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output141_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output142_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output156_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output157_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output158_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output166_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output167_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output171_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output172_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output173_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output177_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output182_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output194_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output196_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output197_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output198_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output199_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output200_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output202_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output208_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1043 ();
endmodule

