* NGSPICE file created from Top_Module_4_ALU.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

.subckt Top_Module_4_ALU ALU_Output[0] ALU_Output[10] ALU_Output[11] ALU_Output[12]
+ ALU_Output[13] ALU_Output[14] ALU_Output[15] ALU_Output[16] ALU_Output[17] ALU_Output[18]
+ ALU_Output[19] ALU_Output[1] ALU_Output[20] ALU_Output[21] ALU_Output[22] ALU_Output[23]
+ ALU_Output[24] ALU_Output[25] ALU_Output[26] ALU_Output[27] ALU_Output[28] ALU_Output[29]
+ ALU_Output[2] ALU_Output[30] ALU_Output[31] ALU_Output[32] ALU_Output[33] ALU_Output[34]
+ ALU_Output[35] ALU_Output[36] ALU_Output[37] ALU_Output[38] ALU_Output[39] ALU_Output[3]
+ ALU_Output[40] ALU_Output[41] ALU_Output[42] ALU_Output[43] ALU_Output[44] ALU_Output[45]
+ ALU_Output[46] ALU_Output[47] ALU_Output[48] ALU_Output[49] ALU_Output[4] ALU_Output[50]
+ ALU_Output[51] ALU_Output[52] ALU_Output[53] ALU_Output[54] ALU_Output[55] ALU_Output[56]
+ ALU_Output[57] ALU_Output[58] ALU_Output[59] ALU_Output[5] ALU_Output[60] ALU_Output[61]
+ ALU_Output[62] ALU_Output[63] ALU_Output[6] ALU_Output[7] ALU_Output[8] ALU_Output[9]
+ Exception[0] Exception[1] Exception[2] Exception[3] Operation[0] Operation[1] Operation[2]
+ Operation[3] Overflow[0] Overflow[1] Overflow[2] Overflow[3] Underflow[0] Underflow[1]
+ Underflow[2] Underflow[3] a_operand[0] a_operand[10] a_operand[11] a_operand[12]
+ a_operand[13] a_operand[14] a_operand[15] a_operand[16] a_operand[17] a_operand[18]
+ a_operand[19] a_operand[1] a_operand[20] a_operand[21] a_operand[22] a_operand[23]
+ a_operand[24] a_operand[25] a_operand[26] a_operand[27] a_operand[28] a_operand[29]
+ a_operand[2] a_operand[30] a_operand[31] a_operand[32] a_operand[33] a_operand[34]
+ a_operand[35] a_operand[36] a_operand[37] a_operand[38] a_operand[39] a_operand[3]
+ a_operand[40] a_operand[41] a_operand[42] a_operand[43] a_operand[44] a_operand[45]
+ a_operand[46] a_operand[47] a_operand[48] a_operand[49] a_operand[4] a_operand[50]
+ a_operand[51] a_operand[52] a_operand[53] a_operand[54] a_operand[55] a_operand[56]
+ a_operand[57] a_operand[58] a_operand[59] a_operand[5] a_operand[60] a_operand[61]
+ a_operand[62] a_operand[63] a_operand[6] a_operand[7] a_operand[8] a_operand[9]
+ b_operand[0] b_operand[10] b_operand[11] b_operand[12] b_operand[13] b_operand[14]
+ b_operand[15] b_operand[16] b_operand[17] b_operand[18] b_operand[19] b_operand[1]
+ b_operand[20] b_operand[21] b_operand[22] b_operand[23] b_operand[24] b_operand[25]
+ b_operand[26] b_operand[27] b_operand[28] b_operand[29] b_operand[2] b_operand[30]
+ b_operand[31] b_operand[32] b_operand[33] b_operand[34] b_operand[35] b_operand[36]
+ b_operand[37] b_operand[38] b_operand[39] b_operand[3] b_operand[40] b_operand[41]
+ b_operand[42] b_operand[43] b_operand[44] b_operand[45] b_operand[46] b_operand[47]
+ b_operand[48] b_operand[49] b_operand[4] b_operand[50] b_operand[51] b_operand[52]
+ b_operand[53] b_operand[54] b_operand[55] b_operand[56] b_operand[57] b_operand[58]
+ b_operand[59] b_operand[5] b_operand[60] b_operand[61] b_operand[62] b_operand[63]
+ b_operand[6] b_operand[7] b_operand[8] b_operand[9] vdd vss
XANTENNA__07383__I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09523__A2 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08326__A3 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05903_ net21 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09671_ _03368_ _03371_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06883_ _00403_ _03955_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06337__A2 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05834_ net79 _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08622_ _01498_ _02231_ _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09304__S _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08553_ _02067_ _02068_ _02142_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05765_ net29 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07504_ _01020_ _01023_ _01024_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_input108_I b_operand[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08484_ _02008_ _02019_ _02081_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05696_ net76 _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07837__A2 _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07435_ _00955_ _00957_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07366_ _00888_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08942__I _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11397__A2 _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09105_ _02753_ _02755_ _02756_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06317_ _03999_ _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07297_ _00819_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08262__A2 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input73_I b_operand[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09036_ _02524_ _02545_ _02680_ _02681_ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06248_ _05459_ _05424_ _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11149__A2 _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06179_ _05392_ net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09762__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _03571_ _03632_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06040__A4 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07293__I _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05806__I _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09514__A2 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09869_ _02429_ _02655_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07525__A1 _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11321__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09013__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10713_ _04365_ _04384_ _04451_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10159__I _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06500__A2 _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ _04363_ _04426_ _04427_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_42_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11388__A2 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10575_ _04351_ _04315_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06264__A1 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10060__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06372__I _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09202__A1 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10899__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11127_ _04893_ _04917_ _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05716__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _04770_ _04776_ _04877_ _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07516__A1 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10009_ _03739_ _03735_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11076__A1 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10823__A1 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08492__A2 _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07220_ _00743_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08762__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07151_ _00668_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09441__A1 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08244__A2 _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06102_ _04086_ _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06255__A1 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ _00538_ _00548_ _00607_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10018__B _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06033_ _04301_ _02997_ _03160_ _04010_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10532__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07984_ _01525_ _01537_ _01538_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_68_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09723_ _03405_ _03413_ _03428_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_47_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06935_ _03683_ _05628_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09654_ _03232_ _00237_ _01189_ _03249_ _03353_ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06866_ _01401_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08605_ _02169_ _02213_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05817_ _02607_ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09585_ _03199_ _03208_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06797_ _00261_ _00303_ _00325_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11067__A1 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08536_ _02117_ _02138_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05748_ _01858_ _01705_ _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10814__A1 _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05679_ _01108_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08467_ _01774_ _02055_ _02056_ _02054_ _02051_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08672__I _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ _00939_ _00940_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08398_ _01934_ _01963_ _01988_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07349_ _00871_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07288__I _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10360_ _04120_ _04121_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09983__A2 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09019_ _02409_ _02563_ _02663_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10291_ _04009_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06706__C1 _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08171__A1 _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10805__A1 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10805__B2 _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06485__A1 _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10281__A2 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10617__I _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10627_ _00675_ _04389_ _04404_ _04409_ net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09423__A1 _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11230__A1 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10033__A2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09974__A2 _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10558_ _04335_ _01417_ _05505_ _03895_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10489_ _04028_ _00232_ _04204_ _04259_ _04260_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05996__B1 _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07737__A1 _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06720_ _00159_ _00163_ _00249_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08757__I _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08162__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06651_ _00169_ _00181_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11049__A1 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06582_ _00083_ _00099_ _00113_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09370_ _02985_ _03043_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08321_ _01904_ _01905_ _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08465__A2 _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08252_ _01829_ _01830_ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07203_ _00651_ _00702_ _00727_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08183_ _01712_ _01755_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09414__A1 _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07134_ _00652_ _00659_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06228__B2 _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07976__A1 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07065_ _00317_ _00580_ _00581_ _00579_ _00577_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_133_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06016_ _01575_ _03030_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09717__A2 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input36_I a_operand[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07967_ _00954_ _00791_ _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09706_ _03406_ _03408_ _03409_ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_74_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06918_ _00358_ _00383_ _00445_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11288__B2 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07898_ _00806_ _01089_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09637_ _03334_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06849_ _02478_ _03356_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07900__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09568_ _03096_ _03109_ _03166_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _02119_ _02120_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09499_ _03174_ _03184_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09653__A1 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08208__A2 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10412_ _04158_ _04163_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_87_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11392_ _05186_ _05199_ _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07967__A1 _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10343_ _04091_ _04093_ _04101_ _04103_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09169__B1 _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09708__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10274_ _03891_ _04028_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07719__A1 _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08931__A3 _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08144__A1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09644__A1 _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11203__A1 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06630__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10082__I _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _02502_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08383__A1 _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07821_ _01361_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07752_ _01239_ _01243_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05904__I _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06703_ _00232_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07683_ _01170_ _01174_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_80_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09422_ _02890_ _02614_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06634_ _00157_ _00164_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09353_ _03022_ _03025_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08438__A2 _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06565_ _00090_ _00093_ _00096_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08304_ _01779_ _01852_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06496_ _05620_ _05622_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09284_ _02903_ _02905_ _02950_ _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_21_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07110__A2 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08235_ _01648_ _01810_ _01811_ _01750_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08166_ _01644_ _01735_ _01736_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07949__A1 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07117_ _00561_ _00565_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08097_ _01588_ _01573_ _01661_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07566__I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07048_ _00573_ _00500_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output142_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08999_ _02471_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06924__A2 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__A1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05814__I _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10961_ _04612_ _04761_ _04771_ _04683_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_43_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06688__B2 _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10484__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10892_ _04605_ _04608_ _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09626__A1 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09626__B2 _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10167__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06860__A1 _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11375_ _05144_ _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10326_ _03823_ _03844_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09157__A3 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10257_ _04006_ _04009_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08365__A1 _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07168__A2 _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08365__B2 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10188_ _03934_ _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06376__B1 _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06915__A2 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08117__A1 _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05724__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08100__I _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07340__A2 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09617__A1 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06350_ _05560_ _02661_ _05302_ _02954_ _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__11424__A1 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10077__I _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06281_ _05462_ _05465_ _05492_ _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_30_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08020_ _00782_ _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08770__I _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06290__I _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07800__B1 _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09971_ _03698_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ _02222_ _02394_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08853_ _02484_ _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07804_ _01330_ _01332_ _01343_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08784_ _02362_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08108__A1 _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05996_ _04539_ _04171_ _04550_ _04215_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07735_ _00762_ _01207_ _01250_ _01268_ net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09856__A1 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07666_ _00899_ _04161_ _01191_ _01193_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10696__B _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09405_ _02998_ _03040_ _03081_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06617_ _00061_ _00120_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09608__A1 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07597_ _01116_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09336_ _02783_ _02386_ _02234_ _03006_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06548_ _00075_ _00079_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09267_ _02924_ _02931_ _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06479_ _05623_ _05631_ _00011_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08680__I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08218_ _00755_ _00931_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09198_ _02782_ _02233_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08149_ _01718_ _00844_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07296__I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08595__A1 _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05809__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11160_ _04897_ _04986_ _04987_ _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10111_ _03848_ _03849_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11091_ _04512_ _03902_ _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10042_ _03690_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07570__A2 _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08855__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10944_ _04748_ _04752_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10875_ _04594_ _04628_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11406__A1 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07086__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06833__A1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11427_ _02152_ _05276_ _05277_ _00735_ net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_125_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05719__I _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11358_ _05146_ _05203_ _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10393__A1 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10309_ _04571_ _04061_ _04062_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11289_ _05115_ _05125_ _05128_ net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08338__A1 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05850_ _02965_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05781_ _02216_ _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07520_ _01039_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08765__I _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08510__A1 _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07451_ _00856_ _00857_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11191__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06402_ _05551_ _05610_ _05611_ _05612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06285__I _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05875__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07382_ _00904_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09121_ _02772_ _02773_ _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06333_ _05543_ _05484_ _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08813__A2 _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06264_ net83 net13 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09052_ _02471_ _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06824__A1 _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08003_ _00814_ _01102_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06195_ _05407_ _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08577__A1 _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10384__A1 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09954_ _03674_ _03679_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08329__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08905_ _02540_ _05497_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09885_ _03573_ _03604_ _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ _02424_ _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10687__A2 _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08767_ _02384_ _02389_ _02252_ _02381_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05979_ _04366_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07718_ _05497_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08675__I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08698_ _02314_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07649_ _01169_ _01175_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06195__I _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10660_ net34 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09319_ _02988_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10591_ _03914_ _04183_ _04123_ _03903_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06815__A1 _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08568__A1 _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11212_ _04950_ _05043_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10375__A1 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11143_ _04886_ _04966_ _04968_ _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09780__A3 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07791__A2 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11074_ _04190_ _04017_ _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput120 b_operand[56] net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput131 b_operand[8] net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_48_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10180__I _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10025_ _03755_ _03756_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10927_ _01430_ _04721_ _04727_ _04097_ _04734_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06319__B _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05857__A2 _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10858_ _04580_ _04631_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_32_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09048__A2 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10789_ _04521_ _04583_ _04584_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06806__A1 _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08559__A1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10366__A1 _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06034__A2 _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07664__I _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06951_ _00364_ _00478_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_79_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05902_ _02564_ _02618_ _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09670_ _03176_ _03369_ _03370_ _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06882_ _03966_ _02085_ _03955_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08621_ _02222_ _02230_ _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05833_ _02780_ _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08552_ _02067_ _02068_ _02142_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05764_ _02031_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05912__I _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07503_ _01001_ _01022_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_63_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08483_ _01993_ _02007_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05695_ _01260_ _01281_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07434_ _00956_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07365_ net129 _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09104_ _02413_ _05586_ _00133_ _02454_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06316_ _05526_ _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07296_ net60 _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08262__A3 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10265__I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09035_ _02589_ _02678_ _02679_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06247_ _05419_ _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input66_I a_operand[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06178_ _05343_ _05391_ _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08014__A3 _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09937_ _03636_ _03638_ _03660_ _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09868_ _03584_ _03586_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_46_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08819_ _02354_ _02408_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09799_ _03413_ _03428_ _03511_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05822__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11085__A2 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ _04365_ _04384_ _04451_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10643_ _04191_ _03868_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10574_ _04351_ _04314_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09169__C _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10175__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06264__A2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10060__A3 _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10348__A1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06016__A2 _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10899__A2 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11126_ _04948_ _04949_ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05775__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11057_ _04772_ _04775_ _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07516__A2 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10008_ _03648_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11076__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10823__A2 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _05344_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09441__A2 _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06101_ _05287_ _05315_ _05316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10085__I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06255__A2 _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07081_ _00524_ _00537_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06032_ _03999_ _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08952__A1 _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07983_ _01333_ _01223_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09722_ _03415_ _03427_ _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06934_ _02269_ _05324_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09653_ _05380_ _03349_ _03350_ _03352_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06865_ _05331_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08180__A2 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08604_ _02175_ _02178_ _02212_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_input120_I b_operand[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05816_ _02596_ _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09584_ _03190_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06738__I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06796_ _00263_ _00302_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08535_ _02122_ _02124_ _02137_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_70_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05747_ _01336_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07062__C _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10814__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08466_ _02046_ _02050_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05678_ _01097_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07417_ _00772_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07691__A1 _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08397_ _01939_ _01962_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07569__I _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07348_ _00870_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10578__A1 _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09432__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07279_ _00796_ _00799_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09018_ _02227_ _02657_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output172_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10290_ _03996_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09196__A1 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05817__I _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08943__A1 _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06706__B1 _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06706__C2 _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08171__A2 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06182__A1 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10805__A2 _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09671__A2 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06485__A2 _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10626_ _04406_ _04407_ _04408_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10569__A1 _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09423__A2 _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11230__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _03884_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10488_ _03917_ _01858_ _04065_ _04615_ _04218_ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__05996__A1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05996__B2 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07737__A2 _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05748__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10741__A1 _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11109_ _04926_ _04928_ _04932_ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06650_ _00172_ _00180_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11049__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06581_ _00105_ _00112_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_45_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__A1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08320_ _00756_ _00770_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09662__A2 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08251_ net71 _00828_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ _00712_ _00721_ _00726_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08182_ _01713_ _01734_ _01754_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07133_ _00654_ _00658_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06228__A2 _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07064_ _00572_ _00576_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10980__A1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06015_ _04495_ _04735_ _04756_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09193__A4 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07966_ _01517_ _01474_ _01518_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09553__B _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09705_ _02286_ _02362_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input29_I a_operand[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ _00359_ _00382_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11288__A2 _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07897_ _00813_ _00829_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09350__A1 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08153__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09636_ _03276_ _03281_ _03333_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_16_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06848_ _00102_ _00367_ _00376_ _00267_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06164__A1 _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07900__A2 _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09567_ _03162_ _03212_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06779_ _00307_ _00308_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09779__I _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08518_ _02032_ _02039_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08683__I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09498_ _03177_ _03180_ _03183_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_70_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10799__A1 _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08456__A3 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08449_ _01986_ _02044_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10411_ _04151_ _04174_ _04175_ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06219__A2 _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11391_ _05237_ _05201_ _05238_ _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10342_ _00992_ _04102_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09169__A1 _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09169__B2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10273_ _03894_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08916__A1 _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06927__B1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08392__A2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07195__A3 _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06942__A3 _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09341__A1 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06155__A1 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09644__A2 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10609_ _04327_ _04331_ _04046_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11203__A2 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10962__A1 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06630__A2 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08907__A1 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08907__B2 _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07820_ _01293_ _01359_ _01360_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08383__A2 _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08768__I _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07751_ _01237_ _01285_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09332__A1 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06702_ _04312_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07682_ _01170_ _01174_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09421_ _03097_ _03099_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06633_ _00159_ _00163_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07894__A1 _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09352_ _02936_ _03024_ _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06564_ _00092_ _00094_ _00095_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_21_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08303_ _01779_ _01852_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07646__A1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09283_ _02913_ _02949_ _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06495_ _01281_ _03705_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08234_ _01747_ _01751_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08165_ _01646_ _01649_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07949__A2 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07116_ _00608_ _00641_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08071__A1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08096_ _01489_ _01500_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10953__A1 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07047_ _00573_ _00500_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10273__I _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10705__A1 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08678__I _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08998_ _02410_ _02640_ _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ _01499_ _01500_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output135_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10960_ _04190_ _04004_ _03859_ _04231_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06137__A1 _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09619_ _03312_ _03315_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_28_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06688__A2 _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10891_ _04605_ _04608_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05830__I _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07637__A1 _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11374_ _05132_ _05218_ _05219_ _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10325_ _03954_ _00950_ _04083_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10256_ _04008_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10187_ _03932_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06376__B2 _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08117__A2 _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06128__A1 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11121__A1 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07876__A1 _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__B2 _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09617__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05740__I _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06280_ _05486_ _05487_ _05491_ _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_30_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10093__I _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07800__A1 _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09970_ _03670_ _03697_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07800__B2 _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08921_ _02397_ _02557_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_112_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08852_ _02248_ _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07616__B _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05915__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07803_ _01340_ _01342_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08783_ _02406_ _02407_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05995_ _02921_ _04539_ _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08108__A2 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ _00816_ _01251_ _01254_ _01255_ _01267_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_37_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11112__A1 _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ _01192_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09404_ _03001_ _03080_ _03039_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06616_ _00036_ _00119_ _00120_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07596_ _01423_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09335_ _02308_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07619__A1 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06547_ _00015_ _00076_ _00078_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10268__I _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input96_I b_operand[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09266_ _02927_ _02930_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07095__A2 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06478_ _05626_ _05630_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08217_ _01787_ _01791_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09197_ _02626_ _02844_ _02855_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06842__A2 _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08148_ net71 _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08595__A2 _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08079_ _01612_ _01641_ _01642_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_1_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10110_ net110 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11090_ _04616_ _04902_ _04911_ _04762_ _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10041_ _02463_ _02406_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__A1 _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10943_ _04700_ _04749_ _04751_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10874_ _04668_ _04676_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10178__I _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07086__A2 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08283__A1 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10090__A1 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06833__A2 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11426_ _05217_ _05275_ _05277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10917__A1 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11357_ _05150_ _05181_ _05201_ _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10308_ _04066_ _00233_ _00414_ _03946_ _04269_ _03836_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11288_ _04842_ _00585_ _05127_ _01255_ _00588_ _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10239_ net41 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07010__A2 _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05780_ net89 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07849__A1 _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08510__A2 _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07450_ _00861_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06401_ _05546_ _05573_ _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_34_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10088__I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07381_ _00903_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09120_ _02352_ _02502_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06332_ _05470_ _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08274__A1 _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08781__I _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09051_ _02645_ _02687_ _02691_ _02698_ net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__10816__I net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06263_ _05471_ _05474_ _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06824__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08002_ _01300_ _01557_ _01558_ _01445_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08026__A1 _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06194_ _02639_ _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09774__A1 _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08577__A2 _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10384__A2 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09953_ _03675_ _03678_ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08904_ _02539_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11333__A1 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09884_ _03591_ _03603_ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07001__A2 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08835_ _02457_ _02460_ _02461_ _02464_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_85_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08766_ _02388_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05978_ _01673_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input11_I a_operand[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09829__A2 _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06760__A1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07717_ _05295_ _01247_ _01248_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08697_ _02312_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07648_ _01170_ _01171_ _01174_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_81_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07579_ _01049_ _00824_ _01050_ _00751_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09318_ _02907_ _02911_ _02987_ _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08265__A1 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10590_ _03903_ _03914_ _04183_ _03950_ _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09249_ _02906_ _02912_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__A1 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11211_ _05011_ _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10375__A2 _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11142_ _04796_ _04967_ _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09780__A4 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09517__A1 _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11073_ _04760_ _04764_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07791__A3 _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput110 b_operand[47] net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput121 b_operand[57] net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput132 b_operand[9] net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10024_ _03685_ _03696_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06751__A1 _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10926_ _04644_ _00966_ _04731_ _04733_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_17_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10857_ _04634_ _04656_ _04657_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10788_ _04519_ _04532_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06806__A2 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08559__A2 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09756__A1 _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11409_ _03852_ _03915_ _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10366__A2 _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09508__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06950_ _00363_ _00476_ _00477_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_98_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11315__A1 _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10118__A2 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I Operation[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05901_ _02737_ _03346_ _03476_ _03520_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_95_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06881_ _00403_ _00408_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08620_ _02229_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05832_ _02769_ _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06742__A1 _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08551_ _02065_ _02147_ _02154_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05763_ _01575_ _02020_ _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07502_ _01021_ _01001_ _01022_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08482_ _02023_ _02041_ _02079_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05694_ _01270_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09692__B1 _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07433_ _00753_ _00768_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07364_ _00886_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09103_ _02754_ _01417_ _05505_ _02452_ _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06315_ _05524_ _05525_ _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09995__A1 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07295_ _00812_ _00817_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09034_ _02678_ _02679_ _02589_ _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06246_ _05456_ _05457_ _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ _05344_ _05373_ _05374_ _05390_ _05391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_2_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input59_I a_operand[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09936_ _02268_ _02540_ _03639_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09867_ net126 _02374_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08686__I _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09291__B _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _02262_ _02271_ _02442_ _02443_ _02446_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_58_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09798_ _03415_ _03427_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08749_ _02370_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10711_ _04454_ _04498_ _04499_ _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10293__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10832__A3 _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10642_ _03887_ _03957_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10045__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10573_ _04294_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10596__A2 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09738__A1 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09202__A3 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08410__A1 _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10191__I _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11125_ _03830_ _03847_ _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08961__A2 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05775__A2 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11056_ _04791_ _04798_ _04874_ _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10007_ _02152_ _03736_ _03737_ _00735_ net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_49_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08477__A1 _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10909_ _04681_ _04715_ _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08229__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09977__A1 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06100_ _03084_ _05314_ _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07080_ _00551_ _00568_ _00605_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06031_ _03008_ _03073_ _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06660__B1 _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08952__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07982_ _00911_ _01375_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06963__A1 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09721_ _03421_ _03426_ _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06933_ _00353_ _00458_ _00460_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09901__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09652_ _03351_ _00232_ _05384_ _02275_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06864_ _05431_ _00392_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08603_ _02127_ _02181_ _02211_ _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_55_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05815_ _02586_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09583_ _03266_ _03275_ _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06795_ _00255_ _00259_ _00323_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input113_I b_operand[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08534_ _02128_ _02136_ _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05746_ _01836_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08465_ _05115_ _02058_ _02061_ net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05677_ _01086_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07416_ _00771_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08396_ _01983_ _01985_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07691__A2 _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07347_ net49 _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09968__A1 _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07278_ _00796_ _00800_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09017_ _02660_ _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06229_ _05439_ _05441_ _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09196__A2 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output165_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08943__A2 _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05757__A2 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09919_ _03633_ _03642_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06706__A1 _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06706__B2 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05833__I _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09120__A2 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07667__C1 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07682__A2 _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10186__I _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10625_ _04406_ _04407_ _04271_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10556_ _04218_ _01073_ _04332_ _01577_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08631__A1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10487_ _03897_ _04257_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05996__A2 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11108_ _05431_ _04931_ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11039_ _04757_ _04802_ _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06580_ _00108_ _00111_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10257__A1 _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08275__B _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08250_ _00784_ net27 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07201_ _00724_ _00725_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08181_ _01737_ _01741_ _01753_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_20_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07132_ _00655_ _00657_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07425__A2 _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08622__A1 _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07063_ _05115_ _00583_ _00589_ net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput200 net200 Exception[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05987__A2 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10980__A2 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06014_ _01477_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09178__A2 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08925__A2 _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10732__A2 _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07965_ _01439_ _01467_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09704_ _02295_ _02350_ _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06916_ _00442_ _00443_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07896_ _01298_ _01441_ _01442_ _01367_ _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10496__A1 _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09350__A2 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09635_ _03303_ _03332_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06847_ _00268_ _02899_ _01531_ _02226_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06778_ _00247_ _00248_ _00306_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09566_ _03218_ _03222_ _03223_ _03217_ _03156_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_83_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08517_ _02034_ _02038_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05729_ _01651_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09497_ _02752_ _03178_ _03181_ _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_23_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08448_ _01989_ _02043_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08861__B2 _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08379_ _01889_ _01891_ _01968_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10410_ _04149_ _04164_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11390_ _05150_ _05181_ _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10341_ _04099_ _04100_ _04071_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09169__A2 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10272_ _03850_ _04025_ _04026_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_79_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08916__A2 _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06927__A1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10723__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06927__B2 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10487__A1 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09341__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07104__A1 _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _04046_ _04327_ _04331_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10539_ _04314_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05738__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10962__A2 _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06091__A1 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08907__A2 _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07750_ _01239_ _01243_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09332__A2 _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06701_ _03900_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07681_ _01169_ _01175_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07343__A1 _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09420_ _03086_ _03098_ _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06632_ _00088_ _00160_ _00162_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08784__I _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09351_ _03023_ _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06563_ _03433_ _05412_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08302_ _01872_ _00421_ _01878_ _01884_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09282_ _02915_ _02948_ _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06494_ _05619_ _05632_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08233_ _00903_ _00888_ _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10650__A1 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08164_ _01646_ _01649_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07115_ _00629_ _00640_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08095_ _01599_ _01659_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07046_ _00435_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09564__B _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input41_I a_operand[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09571__A2 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08997_ _02624_ _02409_ _02378_ _02399_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_76_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07582__A1 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ _00793_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10469__A1 _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06137__A2 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07879_ _00802_ _01349_ _00801_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09618_ _03308_ _03314_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_16_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10890_ _04682_ _04694_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05896__A1 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09549_ _03238_ _05583_ _03239_ _02546_ _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10641__A1 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11373_ _05133_ _05134_ _05205_ _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10944__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10324_ _04066_ _00734_ _04074_ _04388_ _04082_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10255_ _04007_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10186_ _03931_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07573__A1 _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06376__A2 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11121__A2 _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07876__A2 _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09078__A1 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07948__I _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11188__A2 _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09250__A1 _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07800__A2 _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08920_ _02552_ _02554_ _02556_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08851_ _02222_ _02229_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_111_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07802_ _00807_ _04161_ _00584_ _01188_ _01341_ _01193_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_84_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05994_ _02976_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08782_ _02352_ _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07733_ _01258_ _01264_ _01266_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07316__A1 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07664_ _04193_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05931__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09403_ _02999_ _02947_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05878__A1 _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06615_ _00143_ _00145_ _05528_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07595_ _01075_ _01066_ _01116_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09608__A3 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06546_ _05622_ _00077_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09334_ _02308_ _02514_ _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07619__A2 _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10623__A1 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06477_ _00002_ _00009_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09265_ _02925_ _02928_ _02929_ _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_21_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08216_ _01789_ _01790_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input89_I b_operand[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09196_ _02656_ net115 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10284__I _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ net70 _01029_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10926__A2 _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08078_ net6 net91 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08595__A3 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07029_ net29 _03030_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08689__I _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10040_ _03757_ _03773_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08347__A3 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07555__A1 _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06002__I _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10942_ _04600_ _04750_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10862__A1 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10873_ _04671_ _04675_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10614__A1 _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08283__A2 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10090__A2 _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06605__C _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10194__I _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11425_ _05217_ _05275_ _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09232__A1 _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11356_ _05184_ _05200_ _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08586__A3 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09783__A2 _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10307_ _03959_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11287_ _05022_ _05023_ _05033_ _05127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10238_ _03989_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07546__A1 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10169_ _03913_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09932__B _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07849__A2 _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06400_ _05546_ _05573_ _05610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_62_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07380_ net67 _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06331_ _05488_ _05490_ _05541_ _05542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09050_ _02406_ _00950_ _02697_ _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06262_ _05472_ _05473_ _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ _01441_ _01446_ _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06193_ _05364_ _05368_ _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08026__A2 _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06037__A1 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09774__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11030__B2 _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09952_ _03676_ _03677_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08903_ _02504_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09883_ _03594_ _03602_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08834_ _02273_ _02463_ _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08765_ _02387_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05977_ _01596_ _04290_ _04344_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06760__A2 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07716_ _01208_ _01182_ _01246_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_54_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08696_ net56 _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07647_ _01031_ _00859_ _01103_ _01172_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ _01071_ _00752_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09317_ _02328_ _02539_ _02912_ _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_90_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06529_ _05669_ _00035_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09462__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09248_ _02907_ _02911_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_output195_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__A2 _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ _02768_ _02806_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11210_ _04953_ _05010_ _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07776__B2 _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11141_ _03871_ _04235_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09308__I _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11072_ _04765_ _04777_ _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09517__A2 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput100 b_operand[38] net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_88_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11324__A2 _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput111 b_operand[48] net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_103_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput122 b_operand[58] net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10023_ _03680_ _03684_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10189__I _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10925_ _04006_ _01493_ _04732_ _01263_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07700__A1 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10856_ _04566_ _04544_ _04635_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A2 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10787_ _04519_ _04532_ _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11260__A1 _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10063__A2 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06267__B2 _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__A1 _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11408_ _04472_ _05255_ _05257_ _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11339_ _05097_ _05105_ _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09508__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11315__A2 _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05900_ _03498_ _03509_ _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06880_ _00407_ _00313_ _03944_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05831_ _02759_ _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11079__A1 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05762_ _02009_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08550_ _02143_ _02153_ _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07501_ _01019_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10826__A1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05693_ net76 _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08481_ _01991_ _02021_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09692__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07432_ _00740_ _00954_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07363_ _00885_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08247__A2 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09444__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09102_ _02328_ _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06314_ _05509_ _02510_ _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07294_ _00816_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09995__A2 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06245_ _05402_ _05374_ _05428_ _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09033_ _02590_ _02593_ _02604_ _02605_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_11_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06176_ _05375_ _05379_ _05386_ _05389_ _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07758__A1 _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09556__C _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10762__B1 _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09128__I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10762__C2 _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09935_ _03565_ _03644_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06981__A2 _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09866_ net127 _02385_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08183__A1 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08817_ _02444_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09797_ _03489_ _03508_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_46_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08748_ net115 _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09278__A4 _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output208_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08679_ _02288_ _02293_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10710_ _04370_ _04455_ _04452_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10293__A2 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10641_ _04365_ _04384_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09435__A1 _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08238__A2 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11242__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07446__B1 _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10572_ _04318_ _04320_ _04349_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07997__A1 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10450__C1 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08946__B1 _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08410__A2 _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06421__A1 _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11124_ _04944_ _04947_ _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_96_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11055_ _04794_ _04797_ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08174__A1 _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10006_ _03657_ _03652_ _03735_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_76_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08098__B _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10808__A1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08477__A2 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09674__A1 _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06488__A1 _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ _04695_ _04714_ _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10839_ _04555_ _04559_ _04549_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_20_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10036__A2 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07437__B1 _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09977__A2 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07988__A1 _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06030_ _04919_ _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06660__B2 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06412__A1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07981_ _01443_ _01447_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06963__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ _03423_ _03424_ _03425_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06932_ _00298_ _00459_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08787__I _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08165__A1 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09901__A2 _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ _02270_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11427__B _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06863_ _00229_ _00239_ _03922_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07912__A1 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08602_ _02195_ _02204_ _02210_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05814_ _02575_ _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09582_ _03268_ _03274_ _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06794_ _01770_ _02118_ _00260_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08533_ _02131_ _02135_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05745_ _01433_ _01444_ _01195_ _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08468__A2 _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input106_I b_operand[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08464_ _01859_ _00585_ _02060_ _01028_ _00588_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05676_ net12 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07415_ _00930_ _00936_ _00937_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10557__I _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08395_ _01917_ _01984_ _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07346_ _00840_ _00863_ _00868_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07979__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07277_ _00799_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input71_I b_operand[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09016_ _02507_ _02655_ _02568_ _02659_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_124_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06228_ _03509_ _05326_ _05440_ _05330_ _05332_ _05318_ _05441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06159_ _05348_ _05372_ _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06403__A1 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output158_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06954__A2 _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09918_ _03639_ _03641_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08156__A1 _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09849_ _03486_ _03541_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06706__A2 _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07667__B1 _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07667__C2 _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10467__I _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09408__A1 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09959__A2 _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10624_ _04134_ _04038_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10555_ _04331_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06642__A1 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06680__I _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10486_ net36 _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11298__I _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06945__A2 _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11107_ _04834_ _04929_ _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08147__A1 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11038_ _04748_ _04752_ _04855_ _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09647__A1 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10257__A2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07200_ _02107_ _02726_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08180_ _01745_ _01748_ _01752_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07131_ _00653_ _00656_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08622__A2 _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07062_ _00416_ _00585_ _00587_ _05317_ _00588_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput201 net201 Overflow[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06013_ _04495_ _04735_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_133_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07189__A2 _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08925__A3 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07964_ _01439_ _01467_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09703_ _03197_ _03406_ _03315_ _03312_ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06915_ _01760_ _02053_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07895_ _01300_ _01369_ _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09634_ _03307_ _03331_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10496__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06846_ _00278_ _00372_ _00374_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06164__A3 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09565_ _03249_ _03253_ _03255_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06777_ _00247_ _00248_ _00306_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08516_ _02082_ _02116_ _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05728_ _01640_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09496_ net119 net53 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09141__I _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08447_ _02023_ _02041_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08861__A2 _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06872__A1 _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ _01893_ _01896_ _01967_ _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_23_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07329_ _00851_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07596__I _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ _04071_ _04099_ _04100_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10271_ _03848_ _03849_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10184__A1 _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06927__A2 _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08129__A1 _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05844__I _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09877__A1 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10487__A2 _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09629__A1 _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07104__A2 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__B1 _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10607_ _04342_ _04346_ _04387_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10538_ _04302_ _04313_ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10469_ _04232_ _04233_ _04238_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08368__A1 _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10660__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07455__B _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09580__A3 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06700_ _05375_ _00228_ _00229_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07680_ _01176_ _01178_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07343__A2 _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06631_ _00016_ _00161_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ _02285_ net48 _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11427__A1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06562_ _02532_ _05328_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08301_ _01880_ _01881_ _01883_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09281_ _02919_ _02933_ _02947_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06493_ _00010_ _00025_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08232_ _01806_ _01808_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10650__A2 _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08163_ _01721_ _01733_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07114_ _00631_ _00639_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08094_ _01602_ _01658_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07045_ _00508_ _00512_ _00571_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07031__A1 _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08996_ _02613_ _02405_ _02410_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07582__A2 _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input34_I a_operand[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ _01489_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07878_ _00801_ _00910_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07334__A2 _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09617_ net122 _02373_ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06829_ _00343_ _00345_ _00357_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_84_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09548_ _03238_ _02438_ _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05896__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09087__A2 _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ _02292_ _02502_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08834__A2 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05839__I _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11372_ _05133_ _05134_ _05205_ _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10323_ _04080_ _00211_ _04204_ _04081_ _00212_ _03817_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_106_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10254_ net43 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10185_ net97 _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11409__A1 _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10880__A2 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09078__A2 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06836__A1 _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10396__A1 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09002__A2 _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08850_ _04571_ _02480_ _02481_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07801_ _00803_ _00907_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08781_ _02348_ _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05993_ _04485_ _04517_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07732_ _01188_ _01265_ _01189_ _01201_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08513__A1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07663_ _00884_ _00894_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10320__A1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09402_ _02992_ _02996_ _03078_ _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06614_ _00144_ _00140_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10871__A2 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07594_ _00827_ _00880_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09333_ _02924_ _02931_ _03003_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06545_ net21 net79 _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06827__A1 _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09264_ _02319_ _02722_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06476_ _00005_ _00008_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08215_ _01742_ _01744_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09195_ _02785_ _02788_ _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08146_ net72 net16 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08077_ net7 _00764_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07028_ _00553_ _00554_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05802__A2 _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07555__A2 _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output140_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08979_ _02353_ _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08504__A1 _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10941_ _04701_ _04297_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10311__A1 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07858__A3 _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10872_ _04599_ _04672_ _04674_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06818__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10614__A2 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07491__A1 _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11424_ _05220_ _05233_ _05274_ _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11355_ _05186_ _05199_ _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09783__A3 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08991__A1 _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10306_ _04059_ _04062_ _04063_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11286_ _05118_ _05124_ _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10237_ _03987_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10168_ _03912_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _03832_ _00950_ _03834_ _03837_ _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06330_ _05487_ _05491_ _05541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06261_ _05407_ net78 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08000_ _00798_ _01089_ _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06192_ _05350_ _05404_ _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10369__A1 _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06037__A2 _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11030__A2 _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09951_ _02272_ _02655_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08902_ _02536_ _02537_ _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09882_ _03597_ _03601_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_97_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06103__I _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08833_ _02462_ _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10541__A1 _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08764_ _02386_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05976_ _04301_ _04334_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07715_ _01208_ _01182_ _01246_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_66_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08695_ _02310_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07646_ _01090_ _01104_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10844__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07577_ _01048_ _01096_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09316_ _02903_ _02983_ _02984_ _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06528_ _00056_ _00059_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09462__A2 _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ _02367_ _02844_ _02909_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06459_ _05612_ _05639_ _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09178_ _02768_ _02806_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output188_I net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _00757_ _00782_ _01615_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11021__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06579__A3 _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11140_ _04883_ _04888_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11071_ _04875_ _04878_ _04891_ _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput101 b_operand[39] net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput112 b_operand[49] net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10022_ _03752_ _03753_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput123 b_operand[59] net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10924_ _04006_ _04048_ _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07700__A2 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10855_ _04545_ _04546_ _04634_ _04635_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10599__A1 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10786_ _03830_ _03862_ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07464__A1 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06267__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11407_ _03992_ _03890_ _05176_ _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06019__A2 _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11338_ _05099_ _05103_ _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10771__A1 _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11269_ _05092_ _05106_ _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05830_ _02748_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05762__I _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11079__A2 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05761_ _01998_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07500_ _00999_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08480_ _02073_ _02077_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05692_ _01130_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07431_ _00953_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07362_ _00884_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09444__A2 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09101_ _02621_ _01073_ _02752_ _01577_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06313_ _02467_ _03585_ _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07293_ _00815_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09032_ _02590_ _02593_ _02604_ _02605_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_06244_ _05455_ _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07207__A1 _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10843__I _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11003__A2 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06175_ _02683_ _01814_ _05388_ _05389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__A2 _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08955__A1 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05769__A1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10762__A1 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10762__B2 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09934_ _03568_ _03643_ _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09865_ _03580_ _03582_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08183__A2 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09380__A1 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08816_ _02259_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09796_ _03492_ _03507_ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08747_ _02365_ _02367_ _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05959_ _04150_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09132__A1 _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08983__I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ _02292_ _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06497__A2 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07694__A1 _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07629_ _01083_ _01109_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10293__A3 _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10640_ _04360_ _04422_ _04423_ _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09435__A2 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07446__A1 _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ _04317_ _04321_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07446__B2 _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10450__B1 _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10450__C2 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09199__A1 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09319__I _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08946__A1 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05847__I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08946__B2 _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11123_ _04945_ _04946_ _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09763__B _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11054_ _04870_ _04871_ _04872_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10505__A1 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08379__B _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10005_ _03657_ _03652_ _03735_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__A2 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09123__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10808__A2 _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09674__A2 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10907_ _04698_ _04712_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07685__A1 _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06488__A2 _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10838_ _01113_ _04638_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07302__I _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09426__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07437__A1 _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10769_ _04001_ _04168_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07437__B2 _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07988__A2 _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06660__A2 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10744__A1 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06412__A2 _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07980_ _01457_ _01533_ _01534_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06931_ _02357_ _03455_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08165__A2 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09650_ _03147_ _04258_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06862_ _03922_ _00229_ _00239_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06176__A1 _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08601_ _02208_ _02209_ _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07912__A2 _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05813_ net84 _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09581_ _03271_ _03273_ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06793_ _00250_ _00305_ _00321_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_82_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08532_ _02132_ _02134_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05744_ _01814_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08463_ _00939_ _02059_ _01870_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07414_ _00932_ _00935_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08394_ _01915_ _01919_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07212__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07345_ _00864_ _00861_ _00867_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07979__A2 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07276_ _00798_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06100__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09015_ _02657_ _02658_ _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06227_ _03356_ _03444_ _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input64_I a_operand[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06158_ _05346_ _05371_ _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06089_ _02769_ _02009_ _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09917_ _02267_ _02504_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09353__A1 _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09848_ _03481_ _03482_ _03480_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06167__A1 _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05914__A1 _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09779_ _03412_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07667__B2 _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08864__B1 _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10623_ _04046_ _04405_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09758__B _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10554_ _04330_ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08092__A1 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10974__A1 _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06642__A2 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10485_ _04254_ _04255_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08919__A1 _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10726__A1 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11106_ _04812_ _04818_ _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08147__A2 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11037_ _03831_ _03855_ _04753_ _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09895__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07741__B _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11206__A2 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07130_ _02183_ _02715_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10965__A1 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07061_ _00234_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput202 net202 Overflow[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06012_ _04680_ _04702_ _04724_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10717__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08386__A2 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09583__A1 _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07963_ _01468_ _01473_ _01515_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09702_ _02277_ _02615_ _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06914_ _00438_ _00441_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07894_ _00798_ _00750_ _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09633_ _03317_ _03318_ _03330_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_55_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06111__I _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06845_ _00177_ _00373_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09564_ _03249_ _03253_ _03254_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06776_ _00250_ _00305_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_24_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ _02103_ _02115_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05727_ _01629_ _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09495_ _03011_ _03178_ _03179_ _03104_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_24_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08310__A2 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ _02024_ _02027_ _02040_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_51_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06321__A1 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08377_ _01906_ _01965_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06872__A2 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07328_ _00850_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08074__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ _00781_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10270_ _04016_ _04022_ _04024_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output170_I net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09574__A1 _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11381__A1 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10184__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08129__A2 _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07888__A1 _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06560__A1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09629__A2 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06177__B _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__A1 _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__B2 _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10606_ _04348_ _04350_ _04386_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08065__A1 _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10537_ _04305_ _04311_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07812__A1 _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10468_ _03819_ _04237_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08368__A2 _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10399_ _04153_ _04158_ _04163_ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__A1 _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08540__A2 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06630_ net22 net79 _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06551__A1 _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05770__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06561_ _00021_ _00091_ _00092_ _05629_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_45_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ _01859_ _01872_ _04593_ _01882_ _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09096__A3 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09280_ _02935_ _02936_ _02946_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06492_ _00012_ _00024_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08231_ _01788_ _01807_ _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_21_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08162_ _01725_ _01732_ _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07113_ _00634_ _00638_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06067__B1 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08093_ _01604_ _01657_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07044_ _00518_ _00570_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08359__A2 _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05945__I _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10072__B _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08995_ _02636_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07946_ _01429_ _01497_ net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input27_I a_operand[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ _01345_ _01352_ _01405_ _01406_ _01422_ net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_110_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10323__C1 _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09616_ _02295_ _02361_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06828_ _00349_ _00356_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09547_ _03236_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06759_ _00175_ _00287_ _00288_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09478_ _03090_ _03132_ _03161_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08429_ _02022_ _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08047__A1 _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10929__A1 _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11371_ _05131_ _05210_ _05216_ _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10322_ _03953_ _03959_ _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_109_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10253_ _04005_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05855__I _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10184_ _03921_ _03929_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06781__A1 _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06686__I _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07730__B1 _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11409__A2 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09078__A3 _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07089__A2 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06127__S _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07310__I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08589__A2 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09786__A1 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09250__A3 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09538__A1 _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07549__B1 _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06370__B _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05765__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07800_ _01337_ _01338_ _01269_ _00237_ _01339_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08780_ _02378_ _02399_ _02404_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_97_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05992_ _04495_ _04506_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07731_ _05436_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08513__A2 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ _01188_ _04334_ _01189_ _00897_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09401_ _02993_ _02995_ _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_53_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06613_ _02346_ _03759_ _03781_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07593_ _01113_ _01114_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09332_ _02927_ _02930_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06544_ _00014_ _00016_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _02332_ _02615_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06475_ _00003_ _00006_ _00007_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08214_ _01642_ _01788_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09194_ _02790_ _02803_ _02852_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08145_ net5 _00777_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07237__C1 _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09856__B _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08076_ _01559_ _01562_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07027_ _00488_ _00494_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11336__A1 _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08978_ _02613_ _02619_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output133_I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07929_ _01479_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_29_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08504__A2 _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10940_ _04673_ _04703_ _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10311__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10871_ _04524_ _04673_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09465__B1 _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06818__A2 _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06455__B _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07491__A2 _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09768__A1 _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11423_ _05235_ _05236_ _05273_ _05274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_137_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11354_ _05190_ _05198_ _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08440__A1 _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10305_ _04059_ _04062_ _00045_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11285_ _04848_ _05122_ _05123_ _05121_ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10236_ net105 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10167_ net35 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06754__A1 _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10550__A2 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10098_ _03836_ _01825_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07305__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06260_ _03182_ _02802_ _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06191_ _05357_ _05370_ _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09759__B2 _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10369__A2 _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08431__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10615__B _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09950_ _02263_ _02375_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08901_ _02490_ _02525_ _02535_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_124_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09881_ _03598_ _03600_ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08734__A2 _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09931__A1 _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08832_ net62 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09931__B2 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06745__A1 _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10541__A2 _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05975_ _04323_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08763_ _02385_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07714_ _01209_ _01245_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08498__A1 _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input129_I b_operand[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08694_ _02309_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07215__I _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07645_ net69 _00886_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07170__A1 _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07576_ _01095_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10057__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09315_ _02905_ _02950_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09998__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06527_ _00058_ _03759_ _04691_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input94_I b_operand[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06458_ _05612_ _05639_ _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09246_ _02352_ _02584_ _02908_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08670__A1 _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11006__B1 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09177_ _02765_ _02832_ _02833_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_119_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06389_ _02521_ _03607_ _04010_ _05599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ _01604_ _01657_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08422__A1 _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08059_ _01551_ _01555_ _01563_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_122_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10780__A2 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11070_ _04882_ _04890_ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_1_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10021_ _03722_ _03730_ _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput102 b_operand[3] net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput113 b_operand[4] net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput124 b_operand[5] net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06736__A1 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08489__A1 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10923_ _04728_ _01417_ _05590_ _04552_ _04730_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10854_ _04011_ _04653_ _04654_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10048__A1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10486__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10785_ _04577_ _04578_ _04579_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10599__A2 _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07795__I _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11406_ _04394_ _04471_ _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10220__A1 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11337_ _05167_ _05179_ _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10771__A2 _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11268_ _05097_ _05105_ _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10219_ _03947_ _03962_ _03967_ _03968_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07744__B _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11199_ _04026_ _04025_ _04055_ _05030_ _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06727__A1 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05760_ _01987_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05950__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10287__A1 _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05691_ _01238_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10826__A3 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07430_ _00743_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10039__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07361_ net65 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09100_ net118 net54 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09444__A3 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06312_ _05446_ _05454_ _05495_ _05496_ _05523_ net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_07292_ _00814_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09031_ _02649_ _02652_ _02676_ _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06243_ _05405_ _05427_ _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08404__A1 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07207__A2 _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06174_ _02726_ _04150_ _05387_ _03324_ _05337_ _01803_ _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__06415__B1 _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05769__A2 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10762__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09933_ _03645_ _03647_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09904__A1 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09864_ _03418_ _03578_ _03581_ _03516_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10514__A2 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09380__A2 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08815_ _02260_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09795_ _03497_ _03506_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08746_ _02366_ _02363_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05958_ _01716_ _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09132__A2 _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08677_ _02290_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05889_ _03389_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07628_ _01081_ _01110_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07694__A2 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08891__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09160__I _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07559_ _01043_ _01044_ _01078_ net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10570_ _04316_ _04347_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07446__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ _02310_ _00217_ _05332_ _02754_ _02891_ _05512_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10450__B2 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09199__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08946__A2 _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06957__A1 _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _04879_ _04881_ _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11053_ _04759_ _04779_ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06709__A1 _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10004_ _03733_ _03734_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_103_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10906_ _04699_ _04711_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07685__A2 _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10837_ _04569_ _04636_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_32_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10768_ _04047_ _04489_ _04561_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10699_ _04047_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06948__A1 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10744__A2 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06930_ _00350_ _00354_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05773__I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I Operation[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09362__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06861_ _00320_ _00389_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07373__A1 _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06176__A2 _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08600_ _00775_ _00825_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05812_ _02553_ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09580_ _03175_ _03271_ _03272_ _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06792_ _00252_ _00304_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05923__A2 _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08531_ _02130_ _02133_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05743_ _01792_ _01803_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08462_ _01872_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08873__A1 _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07413_ _00932_ _00935_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10680__A1 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08393_ _01910_ _01981_ _01982_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07344_ _00745_ _00769_ _00866_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10432__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07275_ _00797_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10983__A2 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09014_ _02249_ _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06226_ _05434_ _05435_ _03422_ _05437_ _05438_ _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06157_ _05350_ _05357_ _05370_ _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08928__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09050__A1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10735__A2 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input57_I a_operand[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06088_ _05302_ _01542_ _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09916_ _03636_ _03638_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09353__A2 _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09847_ _03470_ _03563_ net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09778_ _03392_ _03398_ _03488_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05914__A2 _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08729_ _02348_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07667__A2 _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08864__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__B2 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08943__B _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10622_ _03896_ _03982_ _03983_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10423__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10553_ _03886_ _04329_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10484_ _04211_ _04217_ _04035_ _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09041__A1 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11105_ _00992_ _04927_ _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09344__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11036_ _04851_ _04852_ _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07355__A1 _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08837__C _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07658__A2 _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10414__A1 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08083__A2 _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05768__I _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07060_ _00586_ _00405_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06011_ _03150_ _04713_ _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput203 net203 Overflow[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09032__A1 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10717__A2 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07594__A1 _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07962_ _01469_ _01472_ _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_96_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09701_ _03317_ _03403_ _03404_ _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06913_ _00439_ _00440_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07893_ _00736_ _00913_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11142__A2 _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09632_ _03328_ _03329_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06844_ net86 _02639_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07897__A2 _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09563_ _05444_ _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06775_ _00252_ _00304_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input111_I b_operand[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08514_ _02105_ _02114_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05726_ _01390_ _01325_ _01618_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09494_ net119 net52 _02373_ net120 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10653__A1 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08445_ _02032_ _02039_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06321__A2 _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08376_ _01908_ _01964_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_104_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10405__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07327_ _00849_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08074__A2 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05678__I _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07258_ _00780_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06209_ _05354_ _05367_ _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07189_ _00629_ _00640_ _00713_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09023__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09574__A2 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output163_I net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07585__A1 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11381__A2 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09326__A2 _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07337__A1 _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06560__A2 _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__A1 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10644__A1 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10605_ _04354_ _04360_ _04385_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08065__A2 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09262__A1 _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09262__B2 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10536_ _04303_ _04308_ _04310_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_109_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10467_ _04235_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09565__A2 _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10398_ _04160_ _04162_ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09317__A2 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11019_ _04015_ _04827_ _03858_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10883__A1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06560_ _03389_ _05407_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06491_ _00013_ _00023_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08230_ net8 _01223_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08161_ _01728_ _01731_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09253__A1 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06067__A1 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11060__A1 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07112_ _00635_ _00637_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08092_ _01606_ _01656_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06067__B2 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07043_ _00520_ _00569_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09556__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08994_ _02354_ _02408_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07945_ _01430_ _01483_ _01485_ _01487_ _01496_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07876_ _00800_ _05644_ _01409_ _05648_ _01421_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_56_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10323__B1 _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10323__C2 _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09615_ _03310_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06827_ _00352_ _00355_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09546_ _02429_ _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06758_ _00103_ _00178_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05709_ net4 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09477_ _03093_ _03131_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_70_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06689_ _00129_ _04290_ _00216_ _00219_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08428_ _01991_ _02021_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08359_ _01718_ _00870_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08047__A2 _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09244__A1 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11370_ _05206_ _05215_ _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10321_ _03941_ _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10252_ _04004_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07558__A1 _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07558__B2 _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10183_ _03925_ _03928_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10562__B1 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06032__I _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06230__A1 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06781__A2 _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05871__I _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07730__A1 _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__B2 _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09078__A4 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07798__I _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06049__A1 _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10519_ _04291_ _04239_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09538__A2 _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07549__A1 _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05991_ _04118_ _02042_ _04182_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06772__A2 _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07730_ _00887_ _00984_ _01262_ _01263_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09710__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07661_ _05519_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09400_ _02989_ _03042_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06612_ _00140_ _00142_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07592_ _01079_ _01080_ _01111_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09331_ _02999_ _02947_ _03001_ _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10608__A1 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06543_ _00012_ _00024_ _00074_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06288__A1 _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09262_ _02779_ _02925_ _02926_ _02859_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06474_ _02489_ _02910_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10348__B _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11408__I0 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08213_ _00789_ _01087_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09226__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09193_ _02662_ _02797_ _02850_ _02851_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_119_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09226__B2 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08144_ _01624_ _01633_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07237__B1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08075_ _01539_ _01636_ _01637_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07026_ _00489_ _00493_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10544__B1 _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06212__A1 _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08977_ _02616_ _02617_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07928_ _01434_ _01478_ _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05691__I _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07859_ _01402_ _01403_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07712__A1 _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10102__I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10870_ net40 net97 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09529_ _03156_ _03217_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08268__A2 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09465__A1 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09465__B2 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07411__I _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09217__A1 _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11422_ _05239_ _05242_ _05272_ _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__11024__A1 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08976__B1 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11353_ _05193_ _05197_ _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08440__A2 _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06451__A1 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10304_ _04061_ _03817_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11284_ _04925_ _05018_ _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11327__A2 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10235_ _03876_ _03885_ _03985_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_106_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06203__A1 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10166_ _03909_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09940__A2 _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07951__A1 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06754__A2 _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10097_ _03825_ _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10838__A1 _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06506__A2 _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07522__S _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08259__A2 _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10999_ _04732_ _04813_ _04726_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_43_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11263__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07321__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11015__A1 _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06190_ _05402_ _05374_ _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06690__A1 _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09759__A2 _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06690__B2 _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05776__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08900_ _02490_ _02535_ _02525_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09880_ _03592_ _03599_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08195__A1 _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ _02304_ _02307_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09931__A2 _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07942__A1 _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08762_ net50 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05974_ _04312_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07713_ _01210_ _01213_ _01244_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_54_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08498__A2 _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08693_ _02308_ _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07644_ _01094_ _01106_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09447__A1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07575_ net124 _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ _02905_ _02950_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10057__A2 _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06526_ _03738_ _05659_ _00057_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09998__A2 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07231__I _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09245_ _02367_ _02844_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06457_ _05665_ _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08670__A2 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11006__A1 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input87_I b_operand[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09176_ _02807_ _02810_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06388_ _02629_ _05597_ _05529_ _03596_ _05598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08127_ _01606_ _01656_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08058_ _01549_ _01617_ _01619_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07009_ _00532_ _00535_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_122_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10020_ _03667_ _03721_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09922__A2 _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput103 b_operand[40] net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput114 b_operand[50] net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_89_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput125 b_operand[60] net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_49_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07933__A1 _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09686__A1 _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10922_ _04722_ _04729_ _04377_ _04730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10853_ _04011_ _04653_ _03254_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10048__A2 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10784_ _04505_ _04534_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11405_ _05249_ _05253_ _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09610__A1 _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08413__A2 _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11336_ _05170_ _05178_ _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10220__A2 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11267_ _05099_ _05103_ _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08177__A1 _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10218_ _03954_ _03960_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_11198_ _05022_ _05029_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07924__A1 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06727__A2 _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10149_ net37 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10287__A2 _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05690_ _01227_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07360_ _00869_ _00879_ _00880_ _00882_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09444__A4 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06311_ _02607_ _05498_ _05501_ _05503_ _05522_ _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07291_ _00813_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09030_ _02669_ _02675_ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06890__I _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06242_ _05449_ _05453_ _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06663__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06173_ _04247_ _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06415__A1 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06415__B2 _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09932_ _03650_ _03653_ _03656_ net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07935__B _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08168__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08610__I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09863_ _02513_ _02255_ _02266_ _02794_ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07915__A1 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08814_ _02265_ _02268_ _02276_ _02440_ _02441_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _03502_ _03505_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08745_ _02356_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09668__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05957_ _04097_ _04129_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08676_ _02289_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05888_ net83 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__A1 _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07627_ _05294_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06351__B1 _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08891__A2 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07558_ _05666_ _01063_ _01067_ _01028_ _01077_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06509_ _00036_ _00041_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07489_ _00945_ _01006_ _01009_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09228_ _02890_ net56 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_139_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10450__A2 _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output193_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09159_ _02814_ _02815_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06406__A1 _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07603__B1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11121_ _04862_ _04880_ _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08159__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11052_ _04801_ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07906__A1 _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10003_ _03658_ _03659_ _03732_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_76_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08331__A1 _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10905_ _04704_ _04707_ _04710_ _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_32_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08882__A2 _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10836_ _04634_ _04635_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10767_ _03998_ _03994_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07437__A3 _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06645__A1 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10698_ _00675_ _04465_ _04477_ _04486_ net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06948__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11319_ _05155_ _05160_ _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06860_ _00322_ _00388_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07373__A2 _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05811_ _02543_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06791_ _00317_ _00319_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08530_ _00781_ _00825_ _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05742_ _01346_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08461_ _02051_ _02057_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08873__A2 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07412_ _00934_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10200__I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06884__A1 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08392_ _01914_ _01933_ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07343_ _00855_ _00865_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09822__A1 _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07274_ net132 _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09013_ _02656_ _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06225_ _03487_ _01227_ _05321_ _05394_ _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06156_ _05358_ _05369_ _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09050__A2 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06087_ _02813_ _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05964__I _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09915_ _03494_ _03637_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09846_ _00425_ _03559_ _03560_ _03562_ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10499__A2 _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09777_ _03395_ _03397_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06989_ _00452_ _00456_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08728_ _02347_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output206_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08659_ net126 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08864__A2 _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10110__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08943__C _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10621_ _04390_ _04392_ _04403_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09813__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10423__A2 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10552_ net37 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10483_ _04253_ _04211_ _04217_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09041__A2 _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05874__I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11104_ _04848_ _04850_ _04925_ _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11035_ _04742_ _04805_ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07355__A2 _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10111__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10819_ _04617_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08607__A2 _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09804__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06618__A1 _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10414__A2 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09280__A2 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06094__A2 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06010_ _03988_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput204 net204 Overflow[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08791__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07961_ _01512_ _01513_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09700_ _03318_ _03328_ _03329_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06912_ _00346_ _00348_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07892_ _01371_ _01389_ _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08543__A1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09631_ _03325_ _03327_ _03322_ _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06843_ _00273_ _00279_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09562_ _02440_ _02556_ _03252_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06774_ _00261_ _00303_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08513_ _02109_ _02113_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05725_ _01607_ _01444_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09493_ net120 net52 _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11026__I _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input104_I b_operand[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08444_ _02034_ _02038_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10653__A2 _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08375_ _01934_ _01963_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05959__I _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07326_ _00848_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07257_ net8 _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06208_ _01270_ _03378_ _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07188_ _00611_ _00627_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07034__A1 _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06139_ _05352_ _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output156_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10105__I _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07337__A2 _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09829_ _03473_ _03544_ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_46_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08837__A2 _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06848__A1 _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05869__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10604_ _04365_ _04384_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09262__A2 _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10535_ _04194_ _04309_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10466_ _04234_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10397_ _03822_ _03927_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08773__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08525__A1 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11018_ _04833_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10883__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07324__I _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06839__A1 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06490_ _00017_ _00020_ _00022_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_33_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05779__I _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08160_ _01723_ _01729_ _01730_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09253__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07111_ _00630_ _00636_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06067__A2 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11060__A2 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08091_ _01616_ _01655_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07042_ _00551_ _00568_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08993_ _02635_ net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10571__A1 _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ _01492_ _01495_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07875_ _01415_ _01419_ _01420_ _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10323__A1 _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10323__B2 _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09614_ _03024_ _03308_ _03309_ _03196_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06826_ _00350_ _00353_ _00354_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_44_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07234__I _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09545_ _03232_ _05589_ _05590_ _03053_ _03234_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_83_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06757_ _00104_ _00178_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05708_ net3 _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09476_ _03158_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06688_ _02247_ _00217_ _00218_ _05330_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08427_ _02008_ _02019_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09229__C1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08358_ net70 _01156_ _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07309_ _00831_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11051__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08289_ _04097_ _01870_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10320_ _02495_ _04078_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10251_ net107 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07409__I _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10182_ _03927_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10562__A1 _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10562__B2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06230__A2 _05429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08507__A1 _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10314__A1 _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10314__B2 _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07730__A2 _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09483__A2 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06049__A2 _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10518_ _04291_ _04239_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08703__I _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10449_ _03905_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08746__A1 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07549__A2 _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05990_ _03063_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07660_ _00812_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06611_ _03770_ _00058_ _00141_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07591_ _05665_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09330_ _02935_ _03000_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06542_ _00013_ _00023_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06893__I _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _02671_ _02310_ _02320_ _02487_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06473_ _02575_ _02759_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08212_ _01737_ _01785_ _01786_ _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09192_ _02798_ _02800_ _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09226__A2 _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08143_ _01635_ _01653_ _01711_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07237__A1 _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07237__B2 _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08074_ _01543_ _01546_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08613__I _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10792__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07025_ _00457_ _00468_ _00466_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06212__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08976_ _02584_ _02542_ _02547_ _02536_ _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input32_I a_operand[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07927_ _01436_ _01476_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_75_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07858_ _01355_ _01358_ _01400_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_56_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07712__A2 _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06809_ _00301_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07789_ _05344_ _01327_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09528_ _03214_ _03216_ _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09465__A2 _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06279__A2 _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ _03056_ _03050_ _03067_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11421_ _05243_ _05246_ _05271_ _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08976__A1 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11352_ _05194_ _05196_ _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10783__A1 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10303_ _04060_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11283_ _04850_ _05121_ _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10234_ _03896_ _03982_ _03983_ _03984_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06203__A2 _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07400__A1 _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _03908_ _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05882__I _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07951__A2 _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05962__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10096_ _03833_ _00734_ _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10838__A2 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08900__A1 _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05714__A1 _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10998_ _04039_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11263__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09208__A2 _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07482__A4 _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06690__A2 _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10526__A1 _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09392__A1 _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08830_ _02458_ _02459_ _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06888__I _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07942__A2 _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08761_ _02383_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05973_ _01629_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09144__A1 _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07712_ _01237_ _01239_ _01243_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_66_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10203__I _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08692_ net120 _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07643_ _01168_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07574_ _01051_ _01054_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ _02835_ _02979_ _02981_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07458__A1 _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06525_ _05650_ _03661_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09244_ _02854_ _02862_ _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06456_ _05294_ _05665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09175_ _02807_ _02810_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11006__A2 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06387_ _05526_ _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08126_ _01599_ _01659_ _01692_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06433__A2 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08057_ _01532_ _01565_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07630__A1 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07008_ _00533_ _00534_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10517__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput104 b_operand[41] net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06197__A1 _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput115 b_operand[51] net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11190__A1 _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput126 b_operand[61] net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08959_ _02480_ _02518_ _02561_ _02598_ _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07697__A1 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10921_ _01792_ _04644_ _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10852_ _04087_ _04651_ _04652_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07449__A1 _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10783_ _04536_ _04574_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10453__B1 _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05877__I _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08949__A1 _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11404_ _05250_ _05251_ _05252_ _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11335_ _05173_ _05177_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07621__A1 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11266_ _05100_ _05102_ _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08177__A2 _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__A1 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10217_ _03963_ _03965_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11197_ _04833_ _04835_ _05027_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10148_ _03890_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09126__A1 _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10079_ _03815_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09677__A2 _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06376__C _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11236__A2 _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06310_ _05508_ _05516_ _05521_ _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07290_ net130 _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06241_ _03531_ _04713_ _05452_ _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06663__A2 _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05787__I _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06172_ _05380_ _05382_ _05385_ _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09601__A2 _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06415__A2 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09931_ _02444_ _00585_ _03655_ _02580_ _00588_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08168__A2 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09862_ _02479_ _02256_ _03578_ _03579_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11172__A1 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08813_ _02274_ _02275_ _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _03500_ _03503_ _03504_ _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_58_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05926__A1 _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09117__A1 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05956_ _04118_ _02042_ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08744_ _02360_ _02364_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08675_ net58 _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05887_ _03367_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08340__A2 _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07626_ _01144_ _01148_ _05663_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06351__A1 _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06351__B2 _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07242__I _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07557_ _01070_ _01076_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06508_ _00040_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07488_ _00854_ _00862_ _01008_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_10_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09227_ net120 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06439_ _02390_ _05505_ _05507_ _05509_ _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09158_ _02749_ _02752_ _02450_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output186_I net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10738__A1 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08109_ _00779_ _01674_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07603__A1 _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10108__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07603__B2 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ _02706_ _02739_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11120_ _04875_ _04942_ _04943_ _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08159__A2 _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _04759_ _04779_ _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11163__A1 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07906__A2 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10002_ _03658_ _03659_ _03732_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07417__I _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08331__A2 _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10904_ _04259_ _04708_ _04709_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_33_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06342__A1 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10835_ _04570_ _04572_ _04632_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08095__A1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10766_ _04042_ _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__A1 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06645__A2 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10697_ _04466_ _04483_ _04484_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09595__A1 _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11318_ _05156_ _05159_ _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08711__I _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11249_ _05080_ _05084_ _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11154__A1 _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09898__A2 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05810_ _02532_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06790_ _00245_ _00307_ _00318_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09542__I _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05741_ _01466_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08460_ _01774_ _02055_ _02056_ _02054_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07411_ _00933_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08391_ _01914_ _01933_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11209__A2 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07342_ _00768_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06636__A2 _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07273_ net68 _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09012_ net53 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ _05436_ _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06155_ _05364_ _05368_ _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06086_ _05300_ _03269_ _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09338__A1 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09914_ _03493_ _03496_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11145__A1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09845_ _00979_ _03561_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _03405_ _03484_ _03485_ _03429_ _03402_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_06988_ _00448_ _00513_ _00514_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05980__I _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08727_ _02345_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05939_ _03900_ _03933_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09510__A1 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08658_ _02265_ _02270_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07609_ _01117_ _01122_ _01132_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08589_ _02103_ _02115_ _02196_ _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08077__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10620_ _04397_ _04398_ _04402_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09813__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10551_ _04326_ _04327_ _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10482_ _04035_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09577__A1 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09627__I _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09329__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11103_ _04848_ _04850_ _04925_ _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11136__A1 _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11034_ _04744_ _04804_ _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06563__A1 _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05890__I _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09501__B2 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06315__A1 _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10111__A2 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10662__A3 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08068__A1 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10818_ _04507_ _04616_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08706__I _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09804__A2 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07815__A1 _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10749_ _04505_ _04534_ _04541_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput205 net205 Underflow[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09537__I _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08791__A2 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07960_ _01436_ _01476_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11127__A1 _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07057__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06911_ _00330_ _00347_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07891_ _01392_ _01398_ _01437_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09630_ _03322_ _03325_ _03327_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09740__A1 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06842_ _00360_ _00365_ _00370_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09272__I _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09561_ _02829_ _02555_ _03251_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06773_ _00263_ _00302_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08512_ _02110_ _02112_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05724_ net3 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09492_ _03165_ _03175_ _03176_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_36_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06306__A1 _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08443_ _02035_ _02037_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08059__A1 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08374_ _01939_ _01962_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08616__I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07520__I _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07325_ net91 _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07256_ _00776_ _00778_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06207_ _05358_ _05369_ _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09559__A1 _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07187_ _00708_ _00709_ _00711_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05975__I _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input62_I a_operand[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06138_ _02889_ _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08231__A1 _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06069_ _04485_ _05158_ _05284_ _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output149_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09828_ _03483_ _03543_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06545__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08300__B _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09759_ _02443_ _00988_ _03467_ _00238_ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10121__I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08298__A1 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09131__B _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10603_ _04368_ _04383_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10534_ _03956_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10465_ net100 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05885__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10396_ _04094_ _04155_ _04159_ _04113_ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_123_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08773__A2 _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11017_ _04023_ _04816_ _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06536__A1 _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10332__A2 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08289__A1 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10096__A1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06839__A2 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06384__C _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09789__A1 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07110_ _02368_ _02489_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ _01620_ _01654_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08461__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07041_ _00552_ _00555_ _00567_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__05795__I _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08213__A1 _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09961__A1 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08992_ _00425_ _02612_ _02630_ _02634_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_88_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07943_ _00921_ _01493_ _00984_ _01337_ _01494_ _01263_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10308__C1 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08516__A2 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09713__A1 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07874_ _01337_ _05517_ _00133_ _01347_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10323__A2 _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _02286_ _02722_ _02486_ _02277_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06825_ _02357_ _05628_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09544_ _03227_ _03233_ _04377_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06756_ _00190_ _00284_ _00285_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05750__A2 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05707_ _01412_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09475_ _03083_ _03089_ _03157_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06687_ _02205_ _03792_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09492__A3 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08426_ _02012_ _02018_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09229__B1 _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09229__C2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08357_ _00784_ _01030_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07308_ _00830_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08288_ _01863_ _01856_ _01867_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07239_ _04919_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10250_ _03864_ _04001_ _04002_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07007__A2 _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10181_ _03926_ _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10116__I _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09704__A1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06518__A1 _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10314__A2 _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06518__B2 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10517_ _04154_ _04232_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06504__I _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10448_ _04216_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08746__A2 _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06757__A1 _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10379_ _04031_ _04141_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10553__A2 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06610_ _02346_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07590_ _01079_ _01080_ _01111_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05732__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06541_ _01760_ _02280_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10608__A3 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09260_ _02308_ _02233_ _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06472_ _05552_ _00003_ _00004_ _05614_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ _01741_ _01753_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09191_ _02730_ _02731_ _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08142_ _01551_ _01555_ _01563_ _01634_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08434__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07237__A2 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06615__S _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10241__A1 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06445__B1 _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08073_ _01543_ _01546_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06996__A1 _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07024_ _00550_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06748__A1 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08975_ _02370_ _02615_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07926_ _01438_ _01475_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input25_I a_operand[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07245__I _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07857_ _01355_ _01358_ _01400_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06808_ _00264_ _00283_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07788_ _01280_ _01248_ _01324_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09527_ _03159_ _03213_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06739_ _00268_ _05352_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09458_ _03056_ _03067_ _03050_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_80_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08409_ _01996_ _02000_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09389_ _03048_ _03064_ _03065_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11420_ _05254_ _05258_ _05270_ _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08425__A1 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10232__A1 _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ _05192_ _05195_ _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08976__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10302_ _03961_ _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11282_ _04934_ _05119_ _05120_ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10233_ _03881_ _03884_ _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10535__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10164_ _03907_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10095_ _03825_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09153__A2 _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07164__A1 _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05714__A2 _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10997_ _04732_ _04726_ _04039_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08714__I _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09613__B1 _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06978__A1 _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10774__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__I _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09916__A1 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08760_ net114 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05972_ _02932_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07711_ _01240_ _01242_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09144__A2 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08691_ _02305_ _02306_ _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07642_ _01155_ _01167_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_80_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06902__A1 _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07573_ _01091_ _01092_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09312_ _02895_ _02980_ _02953_ _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06524_ _02346_ _03770_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09243_ _02327_ _02503_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06455_ _03738_ _05661_ _05663_ _05664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08407__A1 _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08624__I _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09174_ _02827_ _02828_ _02830_ _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06386_ _05588_ _02434_ _05596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10214__A1 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08125_ _01602_ _01658_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09080__A1 _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08056_ _01532_ _01565_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07007_ _00268_ _05407_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10517__A2 _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06197__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput105 b_operand[42] net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07394__A1 _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput116 b_operand[52] net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput127 b_operand[62] net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08958_ _02597_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07909_ _00894_ net49 _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08889_ _02502_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_56_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09686__A3 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10920_ _03855_ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07697__A2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10851_ _04003_ _04265_ _04479_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_71_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07449__A2 _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10782_ _04505_ _04534_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10453__A1 _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10453__B2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11403_ _03862_ _03890_ _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08949__A2 _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__A1 _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10756__A2 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11334_ _05174_ _05176_ _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06054__I _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11265_ _05098_ _05101_ _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05893__I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10216_ _03964_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11196_ _04023_ _04816_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__A1 _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11181__A2 _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10147_ _03888_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09126__A2 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10078_ _03814_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08885__A1 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05699__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10444__A1 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06240_ _04010_ _05451_ _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06171_ _03487_ _04323_ _05384_ _02683_ _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07612__A2 _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09930_ _03654_ _03560_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09365__A2 _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09861_ net128 _02486_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11172__A2 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ _02428_ _02437_ _02439_ _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09792_ _02312_ _02782_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09117__A2 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08743_ _02363_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05955_ _01130_ _04107_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input127_I b_operand[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _02287_ _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09224__B _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08876__A1 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05886_ _03356_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10683__A1 _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07625_ _01144_ _01148_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06887__B1 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07556_ _01072_ _05326_ _01073_ _00832_ _01075_ _05512_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_81_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06139__I _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10435__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06507_ _00038_ _00039_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07487_ _01007_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input92_I b_operand[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05978__I _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09226_ _02306_ _05435_ _02886_ _01123_ _02887_ _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06438_ _05502_ _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_21_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05862__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09157_ _02451_ _02749_ _02752_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__09053__A1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06369_ _05500_ _05514_ _05527_ _05580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__10738__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08108_ _00776_ _00928_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07603__A2 _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08800__A1 _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09088_ _02707_ _02738_ _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_output179_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08039_ _01480_ _01482_ _01570_ _01598_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_116_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11050_ _04867_ _04868_ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11163__A2 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10001_ _03662_ _03664_ _03731_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08867__A1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10903_ _03892_ _04439_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06342__A2 _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10834_ _04573_ _04633_ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10765_ _04493_ _04558_ net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05888__I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07842__A2 _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10696_ _04466_ _04483_ _04271_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09044__A1 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09595__A2 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11317_ _05154_ _05157_ _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11248_ _05081_ _05083_ _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11179_ _04985_ _05008_ _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05740_ _01770_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08858__A1 _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10665__A1 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07410_ net74 _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08390_ _01977_ _01979_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10918__B _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07341_ _00841_ _00843_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08086__A2 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11090__A1 _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07272_ _00791_ _00794_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09011_ _02361_ _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06223_ _01683_ _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10209__I _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06154_ _05354_ _05366_ _05367_ _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_117_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06085_ _01097_ _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09338__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09913_ _03489_ _03634_ _03635_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09844_ _02262_ _03448_ _03442_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06021__A1 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09775_ _03413_ _03428_ _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06987_ _00451_ _00469_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_27_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08726_ _02344_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05938_ _03878_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07253__I _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09510__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08657_ _02268_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05869_ net17 _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07608_ _01126_ _01131_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08588_ _02086_ _02101_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07539_ _01057_ _01058_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08077__A2 _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11081__A1 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10550_ _04255_ _04259_ _04029_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09209_ _02229_ _02315_ _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10119__I net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10481_ _04223_ _04226_ _04251_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06260__A1 _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11102_ _04853_ _04924_ _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11136__A2 _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11033_ _04737_ _04807_ _04849_ _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08001__A2 _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10895__A1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06563__A2 _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09501__A2 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07512__A1 _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10817_ _04614_ _03810_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__A1 _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11072__A1 _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ _04535_ _04536_ _04540_ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10679_ _04395_ _04466_ _04391_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__08722__I _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07579__A1 _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput206 net206 Underflow[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_126_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11288__C _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11127__A2 _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06910_ _00343_ _00436_ _00437_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07890_ _01302_ _01319_ _01391_ _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06841_ _00366_ _00369_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09740__A2 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10699__I _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07751__A1 _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09560_ _02436_ _03243_ _03250_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06772_ _00264_ _00283_ _00301_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08511_ _02104_ _02111_ _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05723_ _01585_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09491_ net56 net116 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06306__A2 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08442_ _02033_ _02036_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_17_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08373_ _01950_ _01961_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07324_ _00846_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07255_ _00777_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06206_ _05406_ _05418_ _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09559__A2 _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07186_ _00529_ _00710_ _00617_ _00615_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08767__B1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06137_ _05136_ _05303_ _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08231__A2 _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07248__I _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input55_I a_operand[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06068_ _02791_ _05180_ _05278_ _05283_ _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09827_ _03486_ _03541_ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06545__A2 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _04571_ _02257_ _02261_ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05753__B1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08709_ _02326_ _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09689_ _03386_ _03391_ _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09495__B2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08807__I _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09247__A1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10602_ _04373_ _04382_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09798__A2 _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05808__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10533_ _04306_ _04307_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10801__A1 _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08470__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06481__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10464_ _03923_ _03957_ _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10395_ _03820_ _03932_ _03951_ _03814_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08222__A2 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09970__A2 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07981__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09373__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10868__A1 _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11016_ _00675_ _04810_ _04825_ _04831_ net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09722__A2 _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10096__A2 _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08717__I _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07040_ _00559_ _00566_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08213__A2 _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09410__A1 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10556__B1 _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ _04919_ _02633_ _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07972__A1 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ _00912_ _00916_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10308__B1 _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10308__C2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ _01416_ _01417_ _01418_ _00796_ _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09612_ net123 _02514_ _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06824_ _03629_ _03237_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09543_ _00213_ _03147_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06755_ _00192_ _00195_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05706_ _01390_ _01401_ _01162_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09474_ _03004_ _03018_ _03088_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06686_ _05279_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10378__B _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08425_ _02014_ _02017_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_24_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09229__A1 _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08356_ _01826_ _01942_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07307_ _00829_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08287_ _01867_ _01863_ _01856_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08452__A2 _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06463__A1 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07238_ _00741_ _01249_ _00748_ _00761_ net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07169_ _05584_ _00693_ _05651_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output161_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ _03920_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07963__A1 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09704__A2 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06518__A2 _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10132__I _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07191__A2 _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__A1 _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08691__A2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11027__A1 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06057__I _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10516_ _03819_ _03888_ _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10447_ _04192_ _04214_ _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09943__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _04140_ _04125_ _04127_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07706__A1 _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06540_ _00069_ _00070_ _00071_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10069__A2 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07351__I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08131__A1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06471_ _05300_ _02423_ _02500_ _01542_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08210_ _01741_ _01753_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06693__A1 _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09190_ _02842_ _02848_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08141_ _01701_ _01709_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08434__A2 _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09631__A1 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06445__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10241__A2 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08072_ _01621_ _01634_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07023_ _00522_ _00549_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10529__B1 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08198__A1 _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09934__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07945__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06748__A2 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08974_ _02614_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07925_ _01439_ _01467_ _01474_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09698__A1 _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07856_ _01362_ _01365_ _01399_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_84_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input18_I a_operand[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06807_ _00334_ _00335_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_28_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07787_ _01280_ _01248_ _01324_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06381__B1 _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11257__A1 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09526_ _03159_ _03213_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_45_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06738_ net88 _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07261__I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08122__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09457_ _03074_ _03137_ _03138_ _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06669_ _00168_ _00199_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_12_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08408_ _01994_ _01997_ _01999_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_51_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11009__B2 _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09388_ _03048_ _03064_ _01139_ _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08339_ _00790_ _01071_ _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09622__A1 _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06436__A1 _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11350_ _04007_ _04195_ _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10232__A2 _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06987__A2 _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10301_ _03836_ _03830_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10127__I _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11281_ _05014_ _05015_ _05013_ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10232_ _03891_ _03895_ _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07936__A1 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06739__A2 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10163_ net99 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07436__I _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09689__A1 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10094_ _03831_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09651__I _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07164__A2 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06911__A2 _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05714__A3 _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10996_ _04738_ _04809_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08113__A1 _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09861__A1 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06675__A1 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__A1 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10759__B1 _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06427__A1 _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06515__I _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06978__A2 _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08730__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05971_ _04279_ _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07710_ _01158_ _01241_ _01222_ _01104_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09144__A3 _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08690_ _02301_ _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08352__A1 _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07641_ _01100_ _01160_ _01166_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_38_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07572_ _00743_ _00821_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08104__A1 _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09311_ _02952_ _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08104__B2 _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06523_ _05662_ _05664_ _00055_ net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07458__A3 _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _02853_ _02875_ _02904_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06454_ _05291_ _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09173_ _02829_ _02455_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09604__A1 _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08407__A2 _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06385_ _05532_ _05533_ _05595_ net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08124_ _01684_ _01686_ _01687_ _01690_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11411__A1 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10214__A2 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09080__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08055_ _01608_ _01615_ _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07006_ _02216_ _05327_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07918__A1 _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput106 b_operand[43] net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07394__A2 _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput117 b_operand[53] net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput128 b_operand[63] net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08957_ _02595_ _02361_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07908_ _01453_ _01454_ _01456_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08888_ _01113_ _02522_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07839_ _01381_ _00829_ _00845_ _00895_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09686__A4 _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10850_ _03864_ _04562_ _04002_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ net121 _02614_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10781_ _04536_ _04574_ _04575_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06657__A1 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08815__I _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11402_ _03989_ _03883_ _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11402__A1 _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__A2 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11333_ _05168_ _05175_ _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09359__B1 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11264_ net42 _04194_ _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A1 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ _03931_ _03939_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09374__A3 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11195_ _03849_ _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08582__A1 _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10146_ _03887_ _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10077_ _03812_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08334__A1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10692__A2 _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10979_ _03898_ _04433_ _03908_ _03892_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08725__I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06170_ _05383_ _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06820__A1 _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09860_ _02255_ _02476_ _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08811_ _02431_ _02438_ _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09791_ _02298_ _02331_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ _02362_ _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05954_ _01749_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08673_ _02286_ _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05885_ net19 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08876__A2 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07624_ _00827_ _00883_ _01008_ _01147_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_81_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10683__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06887__B2 _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07555_ _01074_ _00874_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06506_ _05641_ _05577_ _05605_ _00037_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06639__A1 _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07486_ _00943_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08635__I _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09225_ _02817_ _01227_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06437_ _05645_ _05646_ _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input85_I b_operand[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09156_ _05344_ _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05862__A2 _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06368_ _04442_ _05578_ _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10199__A1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10199__B2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08107_ _01593_ _01594_ _01672_ net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09087_ _02710_ _02736_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_107_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08800__A2 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06299_ _05510_ _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08038_ _01508_ _01595_ _01597_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10000_ _03722_ _03730_ _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09989_ _03703_ _03718_ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10371__A1 _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08316__A1 _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10140__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10902_ _04393_ _04306_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06878__A1 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10833_ _04632_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09816__A1 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10764_ _01430_ _04547_ _04551_ _02495_ _04557_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10695_ _04478_ _04087_ _04482_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06065__I _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05853__A2 _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07055__A1 _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11316_ _04017_ _03938_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11247_ _03872_ _03888_ _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11178_ _04996_ _05007_ _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10362__A1 _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10129_ _03869_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08858__A2 _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06869__A1 _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09807__A1 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06684__B _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07340_ _00841_ _00843_ _00854_ _00862_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08086__A3 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07271_ _00793_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09010_ _02488_ _02509_ _02568_ _02597_ _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_06222_ _01640_ _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06153_ _02769_ _05126_ _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06084_ _05039_ _05049_ _05298_ _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06703__I _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10225__I _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09912_ _03492_ _03507_ _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08546__A1 _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09843_ _03448_ _03442_ _02262_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10353__A1 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09774_ _03413_ _03428_ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06986_ _00451_ _00469_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08725_ net117 _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05937_ _03889_ _03911_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06309__B1 _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__A2 _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ _02267_ _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05868_ _02878_ _03117_ _03160_ _03106_ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07607_ _01068_ _05320_ _00988_ _00825_ _01129_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_54_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ _02182_ _02188_ _02193_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05799_ _02412_ _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07538_ net69 _00871_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06088__A2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07285__A1 _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11081__A2 _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07469_ _00967_ _00734_ _00987_ _00990_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09208_ _02228_ _02314_ _02325_ _02485_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_output191_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10480_ _04241_ _04248_ _04250_ _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_10_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09139_ _02248_ _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_120_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08785__A1 _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11384__A3 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11101_ _04856_ _04923_ _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06260__A2 _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11032_ _04739_ _04740_ _04806_ _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06012__A2 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10895__A2 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07444__I _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07512__A2 _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05899__I _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10816_ net106 _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10747_ _04435_ _04537_ _04538_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_43_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07815__A3 _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10678_ _04044_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09568__A3 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07579__A2 _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__A1 _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput207 net207 Underflow[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10583__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06251__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08528__A1 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06840_ _00367_ _00368_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10886__A2 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07354__I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06771_ _00286_ _00289_ _00300_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_95_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08510_ _01335_ _00806_ _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05722_ _01575_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09490_ net57 net115 _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08700__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08441_ _00789_ _00824_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08372_ _01953_ _01960_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09256__A2 _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07323_ _00845_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11063__A2 _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08464__B1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07254_ net73 _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06205_ _05363_ _05411_ _05417_ _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07185_ _02074_ _02780_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07529__I _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08767__A1 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06136_ _05306_ _05310_ _05349_ _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08767__B2 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06067_ _02845_ _05280_ _05234_ _05282_ _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input48_I a_operand[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10326__A1 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09826_ _03510_ _03540_ _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07264__I _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07742__A2 _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09757_ _02446_ _00414_ _04215_ _02257_ _00235_ _03351_ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_06969_ _00475_ _00496_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05753__B2 _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08708_ _02325_ _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09688_ _03388_ _03390_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08298__A3 _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output204_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _02249_ _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09247__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10601_ _04379_ _04381_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10532_ net33 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10801__A2 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08823__I _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10463_ _03908_ _04231_ _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06481__A2 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10394_ _04154_ _04157_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07981__A2 _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10317__A1 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05992__A1 _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _04813_ _04829_ _04830_ _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07497__A1 _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11293__A2 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11045__A2 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08997__A1 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10484__B _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07349__I _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10556__B2 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08990_ _02613_ _02405_ _02632_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07941_ _04150_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10308__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10308__B2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09174__A1 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10859__A2 _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07872_ _05504_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09611_ _03199_ _03208_ _03306_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06823_ _00194_ _00350_ _00351_ _00297_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_68_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09542_ _02463_ _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06754_ _00192_ _00195_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08908__I _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05705_ _01325_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09473_ _03079_ _03154_ _03155_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06685_ _00210_ _00211_ _00212_ _00048_ _00215_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11284__A2 _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input102_I b_operand[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08424_ _02015_ _02016_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09229__A2 _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ _01824_ _01940_ _01941_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_32_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07306_ _00828_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08286_ _00773_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07237_ _00754_ _01662_ _01738_ _00758_ _00741_ _00760_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_30_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07259__I _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07168_ _03705_ _02607_ _00637_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09401__A2 _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06119_ _05323_ _05333_ _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07099_ _00620_ _00624_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output154_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09809_ _02272_ _02515_ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09468__A2 _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07722__I _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07479__A1 _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11027__A2 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10786__A1 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10515_ _04243_ _04286_ _04287_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10446_ net35 _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10377_ _03935_ _04080_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07954__A2 _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05965__A1 _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05965__B2 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07632__I _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06390__A1 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ _02412_ _05413_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06142__A1 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07890__A1 _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08140_ _01703_ _01708_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08071_ _01624_ _01633_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06445__A2 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07022_ _00538_ _00548_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10529__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10529__B2 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09294__I _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07945__A2 _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08973_ net51 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09147__A1 _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07924_ _01468_ _01473_ _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07855_ _01392_ _01398_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06806_ _01749_ _03856_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07786_ _01323_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06381__A1 _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06381__B2 _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09525_ _03162_ _03212_ _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11257__A2 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06737_ net87 _05213_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09456_ _03074_ _03137_ _04442_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06668_ _00182_ _00198_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08407_ _00933_ _01088_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11009__A2 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09387_ _03060_ _03062_ _02699_ _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06599_ _05504_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05997__I _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08338_ _01813_ _01921_ _01924_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10768__A1 _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09622__A2 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07633__A1 _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08269_ _01795_ _01849_ _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10300_ _03846_ _04056_ _04057_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11280_ _05014_ _05015_ _05013_ _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10231_ _03906_ _03918_ _03980_ _03981_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05946__B _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11193__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10162_ _03901_ _03905_ _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10940__A1 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ _03830_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__I _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10299__B _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10995_ _04807_ _04808_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09861__A2 _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09613__A2 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10759__A1 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10759__B2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07624__A1 _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10429_ _04191_ _04195_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05970_ _01216_ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07640_ _01163_ _01164_ _01165_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07362__I _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07571_ _01053_ _01084_ _01090_ _01013_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10002__B _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08104__A2 _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09310_ _02978_ _02955_ _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06522_ _05666_ _00042_ _00044_ _00047_ _00054_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_62_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09852__A2 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09241_ _02849_ _02876_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06453_ _03738_ _05661_ _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07863__A1 _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09289__I _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09172_ _02447_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06384_ _05577_ _05579_ _05582_ _05317_ _05594_ _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08123_ _00928_ _04161_ _01689_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11411__A2 _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08054_ _01610_ _01614_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07005_ _03651_ _05560_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05929__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10922__A1 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput107 b_operand[44] net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput118 b_operand[54] net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_103_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08956_ _02225_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput129 b_operand[6] net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input30_I a_operand[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07907_ _00903_ net91 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08887_ _02511_ _02517_ _02519_ _02506_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_29_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09540__A1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10686__B1 _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07838_ _01095_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07769_ _00811_ _00765_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09508_ _03114_ _02477_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10780_ _04535_ _04540_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07854__A1 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09439_ _02289_ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06657__A2 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11401_ _03849_ _03941_ _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10138__I _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07606__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11402__A2 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11332_ _03872_ _03879_ _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09359__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11263_ _04007_ _03923_ _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07909__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10214_ _03934_ _03940_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_79_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11194_ _05022_ _05023_ _05024_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10913__A1 _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10145_ _03886_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08582__A2 _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10076_ _03811_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10978_ _04787_ _04790_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_31_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09047__B1 _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08741__I _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07073__A2 _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08022__B2 _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10904__A1 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08573__A2 _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08810_ _02435_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _03499_ _03396_ _03501_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08741_ _02361_ _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05953_ _04086_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08672_ _02285_ _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05884_ _03171_ _03291_ _03313_ _03335_ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__06336__A1 _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07623_ _01008_ _01146_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06887__A2 _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07554_ net49 _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09825__A2 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06505_ _05605_ _00037_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07485_ _00972_ _00867_ _01005_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06639__A2 _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09224_ _00418_ _02311_ _02827_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06436_ _05524_ _05581_ _05596_ _05646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09589__A1 _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06367_ _05534_ _05535_ _05576_ _05578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09155_ _02765_ _02807_ _02810_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10199__A2 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08106_ _01152_ _01660_ _01665_ _01028_ _01671_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08261__A1 _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08651__I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input78_I b_operand[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06298_ _01629_ _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09086_ _02716_ _02735_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08037_ _01512_ _01513_ _01569_ _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11148__A1 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07267__I _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08564__A2 _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09988_ _03709_ _03717_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10371__A2 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08939_ _02547_ _02536_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08316__A2 _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09513__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11320__A1 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10901_ _04216_ _04705_ _04606_ _04706_ _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_44_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10832_ _04576_ _04580_ _04631_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_32_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10763_ _04554_ _04556_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10694_ _04265_ _04479_ _04481_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11315_ _03852_ _03926_ _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08004__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11246_ _04394_ _05076_ _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08555__A2 _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11177_ _04999_ _05005_ _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10362__A2 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10128_ _03868_ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10059_ _03791_ _03793_ _03794_ _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_76_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06318__A1 _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07515__B1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10665__A3 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08736__I _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09807__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10822__B1 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07270_ _00792_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06097__A3 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06221_ _02564_ _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06152_ _05365_ _01987_ _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06083_ _05028_ _05060_ _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09911_ _03508_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09842_ _03555_ _03558_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06557__A1 _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10353__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _03481_ _03482_ _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ _00509_ _00511_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input132_I b_operand[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08724_ _02337_ _02342_ _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05936_ _03900_ _03878_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06309__A1 _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11302__A1 _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08655_ _02266_ _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05867_ _03063_ _03150_ _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07606_ _01879_ _01128_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08586_ _02189_ _02191_ _02192_ _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_05798_ _02401_ _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07537_ _00994_ _01052_ _01056_ _01014_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07285__A2 _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07468_ _00852_ _00988_ _00985_ _00989_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09207_ _02728_ _02798_ _02800_ _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06419_ _05628_ _03193_ _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07399_ _00920_ _00921_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09138_ _02512_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output184_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10041__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09982__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__A2 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09069_ _02653_ _02668_ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11100_ _04858_ _04922_ _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08537__A2 _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09734__A1 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11031_ _04659_ _04720_ _04809_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_77_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10151__I _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10815_ _03998_ _03945_ _04612_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06076__I _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10746_ _04434_ _04436_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10677_ _04413_ _04463_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08225__A1 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10032__A1 _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07579__A3 _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput208 net208 Underflow[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09973__A1 _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10583__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11229_ _03851_ _04307_ _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10335__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07200__A2 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06770_ _00293_ _00296_ _00299_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_48_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10099__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05721_ _01564_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06695__B _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08440_ _00780_ _01071_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08700__A2 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07370__I _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08371_ _01954_ _01959_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07322_ _00844_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08464__A1 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08464__B2 _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10271__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07253_ _00775_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06204_ _05414_ _05415_ _05416_ _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07184_ _00534_ _00621_ _00624_ _00620_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07019__A2 _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06135_ _01749_ _03215_ _05308_ _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09964__A1 _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08767__A2 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10236__I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06066_ _05281_ _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10326__A2 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09825_ _03512_ _03539_ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09756_ _04919_ _03463_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06968_ _00485_ _00495_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_73_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06950__A1 _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05753__A2 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08707_ _02323_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05919_ _03705_ _03716_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ _02940_ _03387_ _02366_ _03287_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06899_ _00322_ _00388_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _02248_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07280__I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08569_ _02170_ _02174_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10600_ _03921_ _04376_ _04380_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08455__A1 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09652__B1 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10531_ net98 _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10462_ _03809_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10146__I _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10393_ _04124_ _04155_ _04156_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_108_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10317__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11014_ _04813_ _04829_ _04271_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07194__A1 _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05703__I _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A1 _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08997__A2 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10729_ _04444_ _04448_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09946__A1 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11202__B1 _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10556__A2 _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07940_ _01490_ _01338_ _00917_ _00237_ _01491_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_141_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10308__A2 _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07365__I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07871_ _05510_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07185__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09610_ _03124_ _03188_ _03304_ _03305_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_95_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06822_ _00295_ _00298_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05735__A2 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09541_ _01118_ _03230_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06753_ _00271_ _00282_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05704_ net1 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09472_ _03153_ _03133_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06684_ _00140_ _00214_ _05245_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08423_ _01334_ _00814_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10492__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10492__B2 _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08354_ net5 net75 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08437__A1 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10244__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07305_ net38 _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06448__B1 _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08285_ _01345_ _01773_ _01854_ _01406_ _01866_ net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_20_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06999__A1 _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07236_ _01825_ _00759_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09937__A1 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07167_ _00600_ _00603_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input60_I a_operand[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06118_ _05325_ _05326_ _05329_ _05330_ _05332_ _02791_ _05333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_07098_ _00622_ _00623_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06049_ _02910_ _05126_ _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output147_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09808_ net125 _02374_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09739_ _02444_ _05589_ _00394_ _03232_ _03446_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07224__B _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__B1 _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10786__A2 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10514_ _04242_ _04246_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_11_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09928__A1 _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10445_ _01423_ _04212_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07939__B1 _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08600__A1 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10376_ _05292_ _04137_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05965__A2 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06142__A2 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08070_ _01627_ _01632_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07642__A2 _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07021_ _00541_ _00547_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10529__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09395__A2 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06602__B1 _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08972_ _02369_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07923_ _01469_ _01472_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07854_ _01393_ _01397_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10701__A2 _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06805_ _00329_ _00333_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ _01284_ _01322_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06381__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09524_ _03168_ _03211_ _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06736_ net89 _01520_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06118__C1 _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09455_ _03135_ _03136_ _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06667_ _00185_ _00197_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06133__A2 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08406_ _00777_ _01030_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08654__I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09386_ _02304_ _02972_ _03061_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07881__A2 _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06598_ _05510_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10217__A1 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08337_ _01751_ _01922_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09083__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07633__A2 _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ _01799_ _01848_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08830__A1 _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ net69 _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08199_ _01767_ _01772_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10230_ _03901_ _03905_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10424__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10161_ _03904_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05947__A2 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10092_ _03827_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08829__I _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08897__A1 _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08649__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06349__I _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10994_ _04739_ _04740_ _04806_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_76_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06124__A2 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05883__A1 _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09074__A1 _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11204__B _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10759__A2 _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07624__A2 _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08821__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09609__B _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ _04194_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _04099_ _04101_ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06060__A1 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08739__I _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08888__A1 _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07570_ _01087_ _01089_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06521_ _00051_ _00053_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09240_ _02902_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06452_ _05658_ _05528_ _05660_ _05661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06520__C1 _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09171_ _02330_ _02415_ _02416_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06383_ _05525_ _05587_ _05593_ _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09604__A3 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08122_ _01879_ _01688_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08812__A1 _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08053_ _01537_ _01611_ _01613_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07004_ _00527_ _00530_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07379__A1 _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08040__A2 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10383__B1 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput108 b_operand[45] net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08955_ _02590_ _02593_ _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput119 b_operand[55] net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07906_ _00796_ _01375_ _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08886_ _02506_ _02511_ _02517_ _02519_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_99_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input23_I a_operand[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10686__A1 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07837_ net129 _00828_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06354__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07768_ _01226_ _01234_ _01304_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09507_ _03113_ _03191_ _03192_ _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06719_ _01770_ _02194_ _00164_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07699_ _01098_ _01228_ _01229_ _01164_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09438_ net59 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05865__A1 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09369_ _02985_ _03043_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11400_ _05161_ _05165_ _05248_ _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07606__A2 _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11331_ _03991_ _03888_ _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10610__A1 _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__I _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09359__A2 _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11262_ _04888_ _05098_ _04972_ _04970_ _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10154__I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10213_ _03954_ _03960_ _03961_ _03946_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11193_ _05022_ _05023_ _00045_ _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10144_ net101 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10075_ _03810_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07463__I _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06345__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10977_ _04750_ _04788_ _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_16_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09295__A1 _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09295__B2 _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05856__A1 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09047__A1 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09047__B2 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09598__A2 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08022__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06033__A1 _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08740_ net52 _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05952_ _04075_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08671_ net122 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05883_ _03324_ _03237_ _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06336__A2 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07622_ _00880_ _01135_ _01145_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07553_ _05506_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06504_ _05640_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07484_ _00967_ _00853_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09223_ _02883_ _02884_ _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10239__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06435_ _05524_ _05581_ _05596_ _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09154_ _02808_ _02738_ _02809_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06366_ _05534_ _05535_ _05576_ _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11396__A2 _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08105_ _01579_ _01238_ _01669_ _01670_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09085_ _02719_ _02734_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08261__A2 _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06297_ _03574_ _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07548__I _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08036_ _01512_ _01513_ _01569_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput90 b_operand[29] net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11148__A2 _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08564__A3 _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09987_ _03711_ _03715_ _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07772__A1 _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06575__A2 _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08938_ _02520_ _02576_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07283__I _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10659__A1 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08869_ _02383_ _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11320__A2 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10900_ _04433_ _04439_ _03913_ _04374_ _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10831_ _04591_ _04630_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10762_ _03990_ _01493_ _00984_ _04400_ _04555_ _01263_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__07827__A2 _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10149__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10693_ _03885_ _04480_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11314_ _04897_ _05154_ _05065_ _05063_ _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11245_ _04903_ _05069_ _05079_ _04991_ _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08004__A2 _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06015__A1 _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10898__A1 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11176_ _05000_ _05004_ _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07763__A1 _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10127_ _03866_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10058_ _02260_ _02377_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07515__A1 _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07515__B2 _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10822__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10822__B2 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08491__A2 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06220_ _05431_ _05432_ _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08752__I _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06151_ _05327_ _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09440__A1 _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06082_ _04843_ _05071_ _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09910_ _03571_ _03632_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10889__A1 _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09841_ _03360_ _03556_ _03557_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06006__B2 _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06557__A2 _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08951__B1 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09772_ _02463_ _02504_ _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06984_ _00444_ _00510_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ _02341_ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05935_ _03856_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07506__A1 _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06309__A2 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input125_I b_operand[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08654_ net63 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05866_ _01292_ _02031_ _03139_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07605_ _01127_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08585_ _00919_ _00807_ _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09259__A1 _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05797_ net86 _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11066__A1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07536_ _00738_ _00835_ _00850_ _00752_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10813__A1 _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07467_ _04204_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input90_I b_operand[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09206_ _02796_ _02865_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06418_ _02694_ _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08662__I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07398_ _00914_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09137_ _02598_ _02659_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06349_ _03433_ _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09431__A1 _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10041__A2 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09068_ _02600_ _02601_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output177_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ _01490_ _01500_ _01577_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11030_ _04842_ _00233_ _04845_ _04604_ _04846_ _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10344__A3 _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08170__A1 _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10814_ _04190_ _03859_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11057__A1 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10745_ _04434_ _04436_ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09670__A1 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10676_ _04461_ _04462_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10032__A2 _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07579__A4 _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11228_ _04895_ _05059_ _05061_ _04986_ _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09725__A2 _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06539__A2 _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07736__A1 _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11159_ net30 net110 _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09489__A1 _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05720_ _01553_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10099__A2 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08161__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06711__A2 _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08370_ _01956_ _01958_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07321_ net27 _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09661__A1 _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08464__A2 _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07252_ _00774_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10271__A2 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06203_ _01097_ _03400_ _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07183_ _00621_ _00703_ _00707_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10559__B1 _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06227__A1 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06134_ _05345_ _05346_ _05347_ _05312_ _04865_ _05071_ _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XANTENNA__09964__A2 _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06065_ _04193_ _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09716__A2 _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10252__I _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _03526_ _03538_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06967_ _00488_ _00494_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09755_ _03459_ _03460_ _02472_ _03462_ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08706_ _02322_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05918_ _03651_ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11287__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09686_ _03120_ _02940_ _03387_ _02358_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__08657__I _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06898_ _00322_ _00388_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08152__A1 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08637_ net112 _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05849_ _02954_ _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08568_ _01413_ _02171_ _02173_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09101__B1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07519_ _00879_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08499_ _02095_ _02097_ _02098_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09652__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09652__B2 _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10530_ _04196_ _04303_ _04304_ _04233_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10461_ _03964_ _04228_ _04229_ _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_108_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ _03940_ _03842_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09707__A2 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11013_ _04014_ _04055_ _04828_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07194__A2 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10728_ _04364_ _04428_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10659_ _03912_ net98 _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06209__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11202__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09946__A2 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11202__B2 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10961__B1 _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07709__A1 _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07870_ _00920_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07185__A2 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ _03553_ _03389_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09540_ _03142_ _03228_ _02436_ _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06752_ _00275_ _00281_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07381__I _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05703_ _01368_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09471_ _03153_ _03133_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06683_ _00213_ _02247_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07488__A3 _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08422_ _01341_ _02010_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06696__A1 _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10492__A2 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08353_ net73 net27 _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07304_ _00822_ _00826_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06448__A1 _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08284_ _01855_ _01857_ _01865_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06448__B2 _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07235_ _00758_ _01890_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07166_ _00686_ _00688_ _00690_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06117_ _05331_ _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07097_ _02324_ _05560_ _05408_ _02237_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input53_I a_operand[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06048_ _02954_ _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07176__A2 _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09807_ net127 _02477_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07999_ _01551_ _01555_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06384__B1 _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09738_ _03440_ _03445_ _05245_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08125__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05804__I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _03288_ _03290_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08428__A2 _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09625__A1 _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__B2 _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09011__I _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07100__A2 _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10513_ _04242_ _04246_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10157__I _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10444_ _04143_ _04210_ _04209_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07939__A1 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07939__B2 _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10375_ _03972_ _04134_ _04135_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08600__A2 _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07466__I _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08364__A1 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07167__A2 _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08116__A1 _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09616__A1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07020_ _00543_ _00546_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08760__I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07376__I _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06602__A1 _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06602__B2 _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08971_ _02609_ _02611_ _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_142_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07922_ _01376_ _01470_ _01471_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09147__A3 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08355__A1 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07853_ _01394_ _01396_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06804_ _00331_ _00332_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07784_ _01286_ _01288_ _01321_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_83_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09523_ _03170_ _03210_ _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06735_ net12 _02140_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06118__B1 _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08658__A2 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06118__C2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09454_ _03076_ _03077_ _03134_ _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09540__B _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06666_ _00186_ _00196_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08405_ _01822_ _01994_ _01995_ _01940_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09385_ _02297_ _02303_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06597_ _02194_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11414__A1 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10217__A2 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08336_ _01334_ _00895_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07995__B _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08267_ _01819_ _01846_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08830__A2 _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07218_ _00739_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08198_ _01137_ _01769_ _01771_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _00670_ _00673_ _00674_ net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08594__A1 _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07286__I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10160_ _03903_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10091_ _03817_ _01662_ _01498_ _03823_ _03828_ _01890_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_59_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10153__A1 _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__A1 _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08649__A2 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10993_ _04739_ _04740_ _04806_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11405__A1 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05883__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09074__A2 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08282__B1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07624__A3 _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08821__A2 _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ _04192_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05709__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10358_ _04115_ _04119_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_98_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10392__A1 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06033__C _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06060__A2 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10289_ _03984_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08888__A2 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06899__A1 _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10695__A2 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06520_ _03716_ _05326_ _00052_ _05330_ _05332_ _05588_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10447__A2 _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09360__B _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08755__I _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06451_ _04702_ _05659_ _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06520__C2 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09170_ _02417_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06382_ _05588_ _05589_ _05590_ _05434_ _05592_ _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08121_ _01666_ _00928_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07076__A1 _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08052_ _01456_ _01612_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07003_ _00525_ _00528_ _00529_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08025__B1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08576__A1 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10383__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10383__B2 _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput109 b_operand[46] net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_130_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08954_ _02559_ _02592_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07905_ net66 _01085_ _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08885_ _02480_ _02518_ _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07000__A1 _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07836_ _01374_ _01376_ _01377_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10686__A2 _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I a_operand[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07767_ _01230_ _01233_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09506_ _03024_ _03115_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06718_ _00154_ _00202_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07839__B1 _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07698_ _00736_ _00888_ _00823_ _01161_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09437_ _03025_ _03116_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06649_ _00175_ _00179_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05865__A2 _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09368_ _02989_ _03042_ _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08319_ _01899_ _01903_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09299_ _02963_ _02966_ _02967_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11330_ _05171_ _05172_ _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11261_ _03991_ _04374_ _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10212_ _03843_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11192_ _04022_ _04929_ _04840_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10374__A1 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10143_ _03881_ _03884_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06042__A2 _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10074_ _03809_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10170__I _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09819__A1 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10429__A2 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10976_ net42 _03948_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09295__A2 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05856__A2 _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09047__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10601__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10904__A3 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06033__A2 _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I a_operand[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05951_ _01618_ _04065_ _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10080__I _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08670_ _02278_ _02283_ _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05882_ _03215_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07621_ _00822_ _00826_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07552_ _01071_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06503_ _05669_ _00035_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07483_ _01004_ net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07836__A3 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _02815_ _02819_ _02827_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06434_ _01727_ _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_107_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07049__A1 _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09153_ _02710_ _02736_ _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06365_ _05538_ _05575_ _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08797__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08104_ _00787_ _00217_ _01667_ _01035_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09084_ _02725_ _02733_ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06296_ _05447_ _05505_ _05507_ _03487_ _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08035_ _01588_ _01592_ _01976_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10255__I _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput80 b_operand[1] net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput91 b_operand[2] net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10356__A1 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09210__A2 _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09986_ _03712_ _03714_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08937_ _02573_ _02574_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10659__A2 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08868_ _04930_ _02474_ _02494_ _02501_ net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07524__A2 _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07819_ _01220_ _01236_ _01296_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_44_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08799_ _02294_ _02425_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08609__B _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10830_ _04592_ _04629_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09277__A2 _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05812__I _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11084__A2 _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10761_ _03990_ _04470_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_40_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10692_ _03881_ _03884_ _03896_ _04274_ _03983_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_40_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07739__I _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11313_ net110 _04309_ _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10165__I _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07460__A1 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11244_ _04990_ _04992_ _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09201__A2 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06015__A2 _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11175_ _05001_ _05003_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10126_ _03865_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07763__A2 _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08960__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10057_ _02273_ _02353_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08712__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07515__A2 _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07279__A1 _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11075__A2 _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10959_ _04689_ _04766_ _04769_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10822__A2 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06150_ _05361_ _05362_ _05363_ _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10586__A1 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06081_ _04865_ _05071_ _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06254__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07203__A1 _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06006__A2 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09840_ _03436_ _03437_ _03435_ _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10889__A2 _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07384__I _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08951__A1 _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09771_ _03479_ _03480_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06983_ _00499_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ _02340_ _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05934_ _03856_ _03878_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08653_ _02264_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05865_ _03019_ _03128_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07604_ _00819_ _01095_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input118_I b_operand[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08584_ _02004_ _02189_ _02190_ _02097_ _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05796_ _02379_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11066__A2 _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07535_ _01051_ _01054_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07466_ _04150_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09205_ _02864_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06417_ _02650_ _05328_ _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07397_ _00919_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input83_I b_operand[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06348_ _02553_ _02009_ _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09136_ _02778_ _02789_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10577__A1 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07442__A1 _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09067_ _02713_ _02714_ _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06279_ _05488_ _05490_ _05491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08018_ _05281_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10329__A1 _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07294__I _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05807__I _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ _03685_ _03696_ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09498__A2 _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10501__A1 _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08170__A2 _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09014__I _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10813_ _04597_ _04610_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_32_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10744_ _03826_ _03991_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09670__A2 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10675_ _04414_ _04416_ _04459_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10280__A3 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09422__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07433__A1 _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06236__A2 _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05995__A1 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09186__A1 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11227_ _04897_ _04987_ _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06322__B _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11158_ net108 net32 _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10109_ _03847_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11089_ _04614_ _04309_ _03810_ _04004_ _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09489__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06172__A1 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11048__A2 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07320_ _00842_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08763__I _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09661__A2 _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ net9 _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06202_ _03258_ _02899_ _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07182_ _00704_ _00705_ _00706_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10559__A1 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10559__B2 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06133_ _05299_ _05311_ _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06227__A2 _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06064_ _05279_ _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05986__A1 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05986__B2 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09823_ _03529_ _03537_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10731__A1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09754_ _02262_ _03461_ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06966_ _00489_ _00493_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08705_ net55 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05917_ _03694_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09685_ _02344_ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06897_ _00244_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07063__B _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08636_ _02245_ _02240_ _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05848_ _02943_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06163__A1 _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08567_ _01271_ _02171_ _01411_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05779_ _02194_ _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09101__A1 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09101__B2 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08673__I _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07518_ _01011_ _01012_ _01038_ net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10798__A1 _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08498_ _00793_ _00886_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09652__A2 _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07663__A1 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07449_ _00762_ _00949_ _00961_ _00971_ net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07289__I _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10460_ _03927_ _04123_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09119_ _02592_ _02770_ _02771_ _02616_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_10391_ _03932_ _03812_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10970__A1 _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__B2 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07238__B _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11012_ _04265_ _04479_ _04827_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08391__A2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06154__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10727_ _04516_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10658_ _04310_ _04438_ _04440_ _04443_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07406__A1 _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11202__A2 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10589_ _03893_ _04295_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10961__A1 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10713__A1 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06820_ _00346_ _00348_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_95_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08758__I _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11269__A2 _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06751_ _00277_ _00280_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_48_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05702_ _01357_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09470_ _03082_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06682_ _01466_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09882__A2 _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08421_ _01830_ _02003_ _02013_ _01946_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_52_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08352_ _01937_ _01938_ _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09634__A2 _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05910__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ _00825_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07645__A1 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08283_ _01685_ _04290_ _01862_ _01864_ _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07234_ _00757_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07165_ _00650_ _00687_ _00689_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06116_ _04236_ _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08070__A1 _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07096_ _00534_ _00621_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__A1 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10263__I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06047_ _05104_ _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input46_I a_operand[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10704__A1 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09806_ _03416_ _03518_ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08668__I _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06384__A1 _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ _01554_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06384__B2 _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09737_ _00213_ _02270_ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06949_ net12 net93 _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09322__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09668_ _02303_ _02349_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09873__A2 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output202_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08619_ _02228_ _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09599_ _03178_ _03181_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10483__A3 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06439__A2 _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10512_ _04278_ _04248_ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_128_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__A1 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10443_ _04143_ _04209_ _04210_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__A2 _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08061__A1 _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10374_ _03972_ _04134_ _04135_ _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08364__A2 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09313__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09616__A2 _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11423__A2 _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10083__I _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06602__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08970_ _02573_ _02610_ _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07921_ _01374_ _01377_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07852_ _01307_ _01395_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10162__A2 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07392__I _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05905__I _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06803_ _00290_ _00292_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput1 Operation[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07783_ _01291_ _01297_ _01320_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09522_ _03186_ _03209_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06734_ _00172_ _00180_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06118__A1 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06118__B2 _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09453_ _03076_ _03077_ _03134_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07866__A1 _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06665_ _00190_ _00192_ _00195_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_input100_I b_operand[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08404_ _01824_ _01941_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09384_ _02304_ _02419_ _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06596_ _00048_ _02335_ _05282_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08335_ _01810_ _01815_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10258__I _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08266_ _01820_ _01845_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07094__A2 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07217_ _00740_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08197_ _00930_ _00946_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08043__A1 _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07148_ _01249_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10925__A1 _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10925__B2 _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08594__A2 _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09791__A1 _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07079_ _00522_ _00549_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output152_I net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10090_ _03825_ _03827_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09543__A1 _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11350__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10153__A2 _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05815__I _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10992_ _04742_ _04805_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_27_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__A2 _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10168__I _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08282__A1 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08282__B2 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06832__A2 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11169__A1 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10426_ net99 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10916__A1 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08585__A2 _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09782__A1 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10357_ _04116_ _04117_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06596__A1 _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10392__A2 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10288_ _04022_ _04039_ _04042_ _04044_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06348__A1 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09298__B1 _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06450_ _02456_ _05598_ _02445_ _05659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06520__B2 _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06381_ _05509_ _04615_ _05591_ _05584_ _05592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08120_ _01666_ _01265_ _01675_ _01123_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08051_ _01333_ _01085_ _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07002_ _03867_ _05352_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08025__A1 _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06291__I _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08025__B2 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08576__A2 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10383__A2 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08953_ _02591_ _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07904_ _01301_ _01370_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08884_ _02516_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11332__A1 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10135__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07835_ _00810_ _00849_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07766_ _01298_ _01299_ _01301_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_37_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09505_ _03024_ _03115_ _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06717_ _00156_ _00201_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07839__A1 _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07839__B2 _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07697_ net129 net16 _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09436_ _03023_ _03113_ _03115_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06648_ _00103_ _00178_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09367_ _02991_ _02998_ _03040_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06579_ _00106_ _00109_ _00110_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__11399__A1 _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09056__A3 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08318_ _01900_ _01902_ _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08681__I _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07067__A2 _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09298_ _02306_ _02822_ _05520_ _02957_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10071__A1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08249_ _00913_ _01102_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07297__I _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11260_ _05094_ _05096_ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10211_ _03959_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_133_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11191_ _03850_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06578__A1 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07775__B1 _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10374__A2 _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10142_ _03883_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 net190 ALU_Output[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09516__A1 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10073_ net31 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06150__B _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09819__A2 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10975_ _04007_ _03841_ _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06502__A1 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08255__A1 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10409_ _04149_ _04164_ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11389_ _05150_ _05181_ _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06569__A1 _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10361__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05950_ _01173_ net2 _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06060__B _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05881_ _02672_ _03302_ _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_39_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ _01143_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06741__A1 _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07551_ _01050_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06502_ _05672_ _00034_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07482_ _00978_ _00982_ _00991_ _01003_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__09691__B1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _02827_ _02815_ _02819_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06433_ _05605_ _05640_ _05642_ _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_61_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08246__A1 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09152_ _02707_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06364_ _05540_ _05542_ _05574_ _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08103_ _01666_ _05191_ _05267_ _01490_ _01668_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09994__A1 _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09083_ _02662_ _02727_ _02732_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06295_ _05506_ _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08034_ _01588_ _01592_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput70 b_operand[10] net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput81 b_operand[20] net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput92 b_operand[30] net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10356__A2 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07221__A2 _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09985_ _03710_ _03713_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_130_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08936_ _02505_ _02236_ _02572_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08867_ _02495_ _02496_ _02499_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07818_ _01220_ _01236_ _01296_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08798_ _02304_ _02419_ _02424_ _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06732__A1 _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07749_ _01213_ _01282_ _01283_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10760_ _04552_ _01338_ _03993_ _05320_ _04553_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09419_ _02322_ _02355_ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10691_ _04051_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08237__A1 _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08788__A2 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10446__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11312_ _05151_ _05152_ _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09737__A1 _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11243_ _05077_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09456__B _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11174_ _04997_ _05002_ _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10125_ net104 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10181__I _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08960__A2 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10056_ _02282_ _02320_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06723__A1 _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08476__A1 _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07279__A2 _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10958_ _04624_ _04768_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10283__A1 _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10889_ _04685_ _04688_ _04693_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08228__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09976__A1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09440__A3 _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06080_ _05294_ _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10305__B _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09770_ _03475_ _03478_ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08951__A2 _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06982_ _00446_ _00498_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06962__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _02339_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05933_ _03867_ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09900__A1 _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08652_ _02263_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05864_ _03030_ _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07603_ _00881_ _00584_ _01120_ _01123_ _01125_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08583_ _02095_ _02098_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05795_ _02368_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09259__A3 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07534_ _00858_ _01052_ _01053_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10274__A1 _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07465_ _00832_ _00983_ _00984_ _00754_ _00986_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09204_ _02799_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06416_ _05481_ _05624_ _05625_ _03280_ _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_10_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ _00918_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10026__A1 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09135_ _02785_ _02788_ _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06347_ _05475_ _05483_ _05557_ _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10266__I _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10577__A2 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input76_I b_operand[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09066_ _02364_ _02383_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06278_ _05409_ _05489_ _05472_ _05367_ _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07442__A2 _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08017_ _01416_ _00126_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09719__A1 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10329__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07575__I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09968_ _03689_ _03695_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06953__A1 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08919_ _02447_ _02555_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09899_ _03619_ _02819_ _03503_ _03620_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_58_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07524__B _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05823__I _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10501__A2 _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10812_ _04598_ _04609_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10743_ _04432_ _04450_ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10674_ _04460_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10017__A1 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__A1 _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05995__A2 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11226_ net110 net31 _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09186__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11157_ _04982_ _04983_ _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06944__A1 _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10740__A2 _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10108_ net46 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11088_ _04773_ _04907_ _04909_ _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10039_ _03758_ _03762_ _03772_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_48_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06172__A2 _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09110__A2 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07250_ _00771_ _00772_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07672__A2 _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06475__A3 _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05683__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ _05412_ _05413_ _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07181_ _02324_ _02553_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10559__A2 _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09875__I _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06132_ _05299_ _05311_ _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07424__A2 _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06063_ _01716_ _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07395__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09822_ _03532_ _03536_ _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06935__A1 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10731__A2 _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09753_ _03440_ _03452_ _02271_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06965_ _00490_ _00492_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input130_I b_operand[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08704_ _02320_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05916_ _03683_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09684_ _02281_ _02392_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08688__A1 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06896_ _00413_ _00415_ _00420_ _00423_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08635_ _02244_ _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05847_ net78 _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08566_ _00920_ _00816_ _02112_ _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05778_ _02183_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09101__A2 _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ _05666_ _01025_ _01027_ _01028_ _01037_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _00914_ _00811_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07448_ _00962_ _00965_ _00970_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07663__A2 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08860__A1 _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07379_ _00812_ _00817_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09118_ _02721_ _02723_ _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output182_I net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10390_ _03819_ _03924_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09049_ _02621_ _05180_ _02695_ _02696_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05977__A2 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A2 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07179__A1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11011_ _04722_ _04651_ _04826_ _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06926__A1 _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08679__A1 _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10726_ _04507_ _04515_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10657_ _03919_ _04441_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08603__A1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__A2 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10588_ _04302_ _04313_ _04367_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10961__A2 _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06090__A1 _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11209_ _04948_ _04949_ _05040_ _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08119__B1 _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06750_ _00273_ _00278_ _00279_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05701_ _01325_ _01346_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06681_ _05331_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08420_ _01945_ _01947_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08351_ _01833_ _01844_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07302_ _00824_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08282_ _00934_ _05280_ _01863_ _05282_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07645__A2 _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08842__A1 _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07233_ _00756_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07164_ _03900_ _05325_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06115_ _05281_ _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06605__B1 _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10401__A1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07802__C1 _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07095_ _02226_ _03367_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10952__A2 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06046_ _01847_ _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input39_I a_operand[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _03515_ _03516_ _03517_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_07997_ _01440_ _01552_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_59_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06948_ net90 net14 _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09736_ _00964_ _03442_ _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10468__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09667_ _03285_ _03301_ _03366_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06879_ _00231_ _03933_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07333__A1 _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08618_ _02227_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08684__I _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09598_ _02309_ _02657_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05895__A1 _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08549_ _02146_ _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07097__B1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10511_ _04226_ _04282_ _04283_ _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10442_ _04033_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10373_ _04031_ _03973_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08061__A2 _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09010__A1 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10459__A1 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08824__A1 _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10709_ _04370_ _04455_ _04452_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_140_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07938__I _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07920_ _01374_ _01377_ _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08769__I _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07851_ _01306_ _01309_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10698__A1 _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11195__I _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07563__A1 _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06802_ _00188_ _00330_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07782_ _01302_ _01319_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput2 Operation[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09521_ _03190_ _03199_ _03208_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06733_ _00182_ _00198_ _00262_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06118__A2 _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09452_ _03079_ _03082_ _03133_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06664_ _05440_ _00193_ _00194_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07866__A2 _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08403_ _00772_ _00749_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10870__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09383_ _03049_ _03051_ _03058_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06595_ _05650_ _00126_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08334_ _01915_ _01919_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08265_ _01833_ _01844_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07216_ _00739_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08196_ _01674_ _01768_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ _00671_ _00672_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08043__A2 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10925__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09791__A2 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07078_ _00600_ _00603_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06029_ _01488_ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09543__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10689__A1 _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output145_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10689__B2 _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10223__B _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11350__A2 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09719_ _02220_ _02263_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10991_ _04744_ _04804_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10310__B1 _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05831__I _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10449__I _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10861__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09459__B _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08282__A2 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11169__A2 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10425_ _04190_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09231__A1 _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09231__B2 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10916__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10356_ _03826_ _03941_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09782__A2 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07793__A1 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10287_ _03869_ _03874_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06348__A2 _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07545__A1 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11341__A2 _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09298__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07442__B _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05741__I _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10852__A1 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06520__A2 _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06380_ _01868_ _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10604__A1 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _01525_ _01538_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07001_ _02140_ _02748_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10094__I _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10368__B1 _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06036__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09773__A2 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08981__B1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08952_ _02359_ _02487_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05916__I _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07903_ _01378_ _01387_ _01450_ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08883_ _02483_ _02488_ _02516_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__07536__A1 _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11332__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07834_ _00804_ _01375_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07765_ _01214_ _01300_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06716_ _00149_ _00204_ _00245_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11096__A1 _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09504_ _03118_ _03187_ _03189_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07696_ _01221_ _01225_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07839__A2 _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09435_ _02219_ _03114_ _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06647_ _00173_ _00176_ _00177_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_24_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09366_ _03002_ _03039_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06578_ _02489_ _02759_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08317_ _01806_ _01808_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09297_ _02964_ _05511_ _01418_ _02303_ _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06275__A1 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08248_ _01822_ _01823_ _01826_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10071__A2 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08179_ _01747_ _01750_ _01751_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10210_ _03958_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11020__A1 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11190_ _01113_ _05020_ _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07775__A1 _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06578__A2 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07775__B2 _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10141_ _03882_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput180 net180 ALU_Output[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05826__I _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput191 net191 ALU_Output[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09516__A2 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10072_ _03807_ _03808_ _00674_ net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10974_ _04688_ _04784_ _04785_ _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10179__I _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__I _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08255__A2 _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06266__A1 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06266__B2 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10408_ _04033_ _04172_ _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11011__A1 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11388_ _04728_ _03910_ _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07766__A1 _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06569__A2 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10339_ _04095_ _04098_ _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05736__I _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11314__A2 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05880_ _02726_ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08191__A1 _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07550_ _01068_ _05435_ _00876_ _05437_ _01069_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_53_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06501_ _05675_ _00033_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10825__A1 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10089__I _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07481_ _00992_ _01001_ _01002_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09691__A1 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09691__B2 _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09220_ _02835_ _02881_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06432_ _05641_ _05577_ _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09151_ _02766_ _02768_ _02806_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06363_ _05546_ _05551_ _05573_ _05574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08246__A2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09443__A1 _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07398__I _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08102_ _00395_ _01667_ _01586_ _00397_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09082_ _02728_ _02730_ _02731_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06294_ _04247_ _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08033_ _01589_ _01591_ _00974_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput60 a_operand[5] net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput71 b_operand[11] net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput82 b_operand[21] net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput93 b_operand[31] net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_1_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07757__A1 _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10552__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09984_ _02290_ _02783_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08935_ _02505_ _02236_ _02572_ _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_57_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08866_ _02497_ _02498_ _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input21_I a_operand[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07861__I _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07817_ _01288_ _01356_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08797_ _02421_ _02422_ _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06732__A2 _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07748_ _01210_ _01244_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07679_ _01154_ _01179_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08692__I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09418_ _02937_ _02371_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10292__A2 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10690_ _03885_ _03985_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__A2 _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _02244_ _02288_ _02305_ _02380_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_138_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11241__A1 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10044__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11311_ _05067_ _05073_ _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11242_ _04913_ _05076_ _05003_ _05001_ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09737__A2 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10462__I _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11173_ net103 net37 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10124_ _03860_ _03863_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10055_ _03615_ _03775_ _03708_ _03704_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_76_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08173__A1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10807__A1 _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10807__B2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10957_ _03865_ net34 _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10283__A2 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10888_ _04617_ _04692_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_129_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09425__A1 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__A2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07987__B2 _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08551__B _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10372__I _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06411__A1 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06981_ _00442_ _00443_ _00507_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06962__A2 _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ _02338_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05932_ net92 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08777__I _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08164__A1 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08651_ net127 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05863_ _03008_ _03073_ _03106_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07602_ _01068_ _05169_ _01124_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08582_ _00786_ _00886_ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05794_ _02357_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07533_ _00830_ _00766_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09664__A1 _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06478__A1 _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ _05202_ _00985_ _00860_ _04377_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10274__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09203_ _02854_ _02862_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06415_ _02704_ _02759_ _02910_ _03400_ _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09416__A1 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08219__A2 _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07395_ net6 _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09134_ _02770_ _02786_ _02787_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06346_ _05479_ _05482_ _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10026__A2 _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09967__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09065_ _02711_ _02712_ _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06277_ _03084_ _05410_ _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08016_ _01572_ _01573_ _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input69_I b_operand[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09719__A2 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06650__A1 _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09967_ _03690_ _03693_ _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_77_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07805__B _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08687__I _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08918_ _02470_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09898_ _03500_ _03504_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08849_ _02475_ _02238_ _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09104__B1 _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10811_ _04601_ _04605_ _04608_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06000__I _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06469__A1 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07666__B1 _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10742_ _04518_ _04533_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10673_ _04414_ _04416_ _04459_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10017__A2 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07969__A1 _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08630__A2 _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06641__A1 _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10406__B _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11225_ _04989_ _04993_ _05057_ _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10192__I _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08394__A1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11156_ _04906_ _04916_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10107_ _03839_ _03844_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10920__I _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11087_ _04690_ _04908_ _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08146__A1 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10038_ _03763_ _03768_ _03771_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_64_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09894__A1 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__A2 _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06200_ _01520_ _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11205__A1 _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09949__A2 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ _03867_ _03204_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06131_ _05297_ _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08621__A2 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06062_ _03324_ _05191_ _03095_ _05256_ _05267_ _04301_ _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09821_ _03533_ _03535_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06935__A2 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09752_ _02271_ _02442_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06964_ _00486_ _00491_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_86_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08137__A1 _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08703_ _02319_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05915_ net23 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09683_ _03311_ _03316_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06895_ _00421_ _00422_ _00417_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08688__A2 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input123_I b_operand[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05846_ _02921_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08634_ _02220_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08565_ _02073_ _02077_ _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05777_ _02172_ _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07516_ _00832_ _04290_ _01034_ _01036_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08496_ _00785_ _00820_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07447_ _00754_ _00966_ _00963_ _04388_ _00969_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_50_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__A2 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06871__A1 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07378_ _00827_ _00883_ _00897_ _00900_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06871__B2 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06329_ _05486_ _05539_ _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09117_ _02345_ _02722_ _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09048_ _02581_ _01410_ _02637_ _04593_ _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_output175_I net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11010_ _04012_ _04048_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07179__A2 _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10183__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06926__A2 _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05834__I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09628__A1 _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08300__A1 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__I _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10725_ _04510_ _04514_ _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_41_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08851__A2 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08880__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10656_ net34 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11199__B1 _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10587_ _04305_ _04311_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06090__A2 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11208_ _04944_ _04947_ _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_122_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11139_ _04959_ _04964_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08119__A1 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09867__A1 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05700_ _01173_ _01336_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10477__A2 _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06680_ _04312_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08350_ _01821_ _01935_ _01936_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11426__A1 _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09095__A2 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07301_ _00823_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10097__I _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08281_ _01685_ _00934_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07232_ _00755_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07163_ _00563_ _00687_ _00657_ _00655_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06605__A1 _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06114_ _05327_ _05328_ _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10401__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07802__B1 _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07094_ _03651_ _02543_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06605__B2 _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07802__C2 _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06045_ _05071_ _05082_ _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08358__A1 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ _02512_ net64 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07030__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07996_ _00792_ _00750_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09735_ _03344_ _03349_ _03440_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06947_ _00473_ _00474_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10468__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09666_ _03286_ _03300_ _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06878_ _04097_ _00405_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08530__A1 _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08617_ _02225_ _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05829_ net15 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09597_ _03288_ _03290_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11417__A1 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08548_ _00951_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07097__A1 _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07097__B2 _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08479_ _02075_ _02076_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10510_ _04223_ _04251_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06844__A1 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10441_ _03930_ _04141_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05829__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10372_ _04027_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09010__A2 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10459__A2 _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08875__I _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08521__A1 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07088__A1 _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08824__A2 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06835__A1 _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10708_ _04421_ _04494_ _04496_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10639_ _04354_ _04385_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_6_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09001__A2 _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10380__I _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07850_ _01305_ _01318_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10698__A2 _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07563__A2 _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06801_ _02269_ _02802_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07781_ _01305_ _01318_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 Operation[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09520_ _03126_ _03200_ _03207_ _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06732_ _00101_ _00104_ _00112_ _00181_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_36_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09451_ _03090_ _03132_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06663_ _02532_ _05412_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08402_ _01943_ _01948_ _01992_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10870__A2 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09382_ _03055_ _03057_ _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06594_ _05387_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08333_ _01917_ _01918_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_32_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08264_ _01838_ _01843_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10555__I _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07215_ _00738_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08195_ _01587_ _01589_ _00779_ _00788_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08579__A1 _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07146_ _00592_ _00669_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07077_ _00601_ _00602_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input51_I a_operand[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06028_ _04528_ _04560_ _04669_ _04898_ net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10689__A2 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07979_ _01460_ _01462_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output138_I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09718_ _02429_ _02515_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08695__I _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10990_ _04754_ _04803_ _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09649_ _02274_ _03232_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10310__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10310__B2 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10861__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09059__A2 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06817__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10465__I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07490__A1 _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10424_ net30 _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10377__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09231__A2 _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10355_ _03821_ _03953_ _03843_ _03815_ _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_83_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06596__A3 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08990__A1 _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10286_ _04040_ _04041_ _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09298__A2 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10301__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07014__I _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07481__A1 _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07000_ _00361_ _00525_ _00526_ _00476_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_116_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09222__A2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10368__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10368__B2 _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07784__A2 _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08981__A1 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08981__B2 _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08951_ _02223_ _02360_ _02584_ _02236_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07902_ _01383_ _01386_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08882_ _02513_ _02515_ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07833_ net80 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10540__A1 _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07764_ _00805_ _00749_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05932__I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09503_ _03027_ _03029_ _03188_ _03123_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_71_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06715_ _00152_ _00203_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11096__A2 _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07695_ _01222_ _01224_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ net123 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06646_ net85 _03182_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06511__A3 _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09365_ _03020_ _03021_ _03038_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_40_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06577_ _02586_ _05365_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08316_ _01788_ _01807_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input99_I b_operand[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09296_ _02293_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10285__I _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06275__A2 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08247_ _01714_ _01824_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07472__A1 _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08178_ _00904_ _01381_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11020__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _02107_ _05325_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10140_ net39 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07775__A2 _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput170 net170 ALU_Output[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput181 net181 ALU_Output[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput192 net192 ALU_Output[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10071_ _03742_ _03806_ _05295_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09516__A3 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05842__I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11087__A2 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10973_ _04617_ _04692_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05998__B _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10598__A1 _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10598__B2 _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06018__A2 _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10407_ _03979_ _04167_ _04168_ _04170_ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_11387_ _05193_ _05197_ _05198_ _05190_ _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10338_ _04095_ _04098_ _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10770__A1 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10269_ _04023_ _04020_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08191__A2 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09140__A1 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06500_ _00001_ _00026_ _00032_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_46_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07480_ _00999_ _01000_ _00958_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10825__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09691__A2 _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ _05538_ _05575_ _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_21_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06362_ _05556_ _05572_ _05573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09150_ _02774_ _02805_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10589__A1 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09443__A2 _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08101_ _01584_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09081_ _02508_ _02341_ _02409_ _02666_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06293_ _05504_ _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08032_ _01501_ _01590_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput50 a_operand[50] net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput61 a_operand[60] net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_128_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput72 b_operand[12] net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_116_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput83 b_operand[22] net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput94 b_operand[32] net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_143_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07757__A2 _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09983_ _02281_ _02334_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__A1 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08934_ _02559_ _02571_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08865_ _02224_ _00235_ _02480_ _00989_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08182__A2 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07816_ _01286_ _01321_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06193__A1 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08796_ _02420_ _02293_ _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input14_I a_operand[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07747_ _01210_ _01244_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09131__A1 _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08973__I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07678_ _01201_ _01206_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_13_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09417_ _03013_ _03017_ _03094_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06496__A2 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06629_ _00077_ _00089_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09348_ _02936_ _02946_ _02945_ _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11241__A2 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09279_ _02939_ _02941_ _02944_ _02872_ _02945_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_32_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11310_ _05062_ _05066_ _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11241_ _03866_ _04329_ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05837__I _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11172_ _03882_ _03887_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10123_ _03862_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08960__A4 _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10054_ _03787_ _03788_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10504__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A2 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09122__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10956_ _04686_ _04690_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10887_ _04686_ _04689_ _04690_ _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09425__A2 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05998__A1 _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08936__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06411__A2 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06980_ _00438_ _00441_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I a_operand[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05931_ net28 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08279__B _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09361__A1 _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08164__A2 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08650_ _02257_ _02261_ _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06175__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05862_ _03084_ _03095_ _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_27_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07601_ _00887_ _04323_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08581_ _02184_ _02185_ _02187_ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_82_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05793_ net22 _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07532_ _00834_ _00751_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09664__A2 _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07463_ _00859_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09202_ _02784_ _02857_ _02861_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06414_ _03389_ _05223_ _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ _00912_ _00916_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09416__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09133_ _02366_ _02375_ _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06345_ _05552_ _05553_ _05555_ _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_120_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__A2 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06276_ _05406_ _05418_ _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09064_ _02670_ _02674_ _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10982__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08015_ _01494_ _01486_ _01502_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08927__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09966_ _03686_ _03691_ _03692_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_77_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08917_ _02525_ _02528_ _02398_ _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09897_ _03006_ _02314_ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09352__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08848_ _02479_ _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08779_ _02400_ _02403_ _02397_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_73_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09104__A1 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10810_ _04603_ _04606_ _04607_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09104__B2 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10741_ _04519_ _04521_ _04532_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07666__A1 _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06469__A2 _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07666__B2 _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10672_ _04421_ _04424_ _04458_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09748__B _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11224_ _04899_ _04988_ _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10725__A1 _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11155_ _04894_ _04980_ _04981_ _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08878__I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10106_ _03843_ _03815_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11086_ net104 net35 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08146__A2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09343__A1 _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10489__B1 _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10037_ _03599_ _03763_ _03769_ _03691_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_48_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10648__I _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10939_ _04698_ _04712_ _04747_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06130_ _01847_ _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08082__A1 _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06061_ _04247_ _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10716__A1 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09820_ _03527_ _03534_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _02446_ _02443_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06963_ net85 net20 _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08137__A2 _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08702_ _02318_ _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05914_ _03629_ _03661_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09682_ _03292_ _03382_ _03383_ _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06148__A1 _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06894_ _03966_ _05380_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09885__A2 _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _02224_ _01249_ _02232_ _02243_ net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05845_ _02910_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07896__A1 _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input116_I b_operand[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08564_ _02164_ _02166_ _02168_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_54_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05776_ net25 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07515_ _00837_ _00217_ _01031_ _01035_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08495_ _02089_ _02093_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07446_ _00967_ _04637_ _00968_ _00741_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07377_ _00898_ _00899_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06871__A2 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input81_I b_operand[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09116_ _02716_ _02735_ _02767_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06328_ _05487_ _05491_ _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08073__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10955__A1 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07820__A1 _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09047_ _02413_ _04637_ _02692_ _02693_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06259_ _03367_ _01987_ _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09948__I0 _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output168_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08376__A2 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08698__I _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10183__A2 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09949_ _03236_ _02351_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09325__A1 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05850__I _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09628__A2 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10724_ _04508_ _04511_ _04513_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06311__A1 _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06311__B2 _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10655_ _04439_ _03938_ _04375_ _03898_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10586_ _04361_ _04362_ _04364_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09261__B1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10946__A1 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08603__A3 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09800__A2 _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07811__A1 _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11207_ _05019_ _05021_ _05025_ _05038_ net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11138_ _04961_ _04963_ _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_122_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08119__A2 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11069_ _04885_ _04889_ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09867__A2 _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10477__A3 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11426__A2 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07300_ net124 _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08280_ _01859_ _00130_ _00212_ _01666_ _01861_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07231_ _00744_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09388__B _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07162_ _02183_ _03509_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10937__A1 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06113_ net81 _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07802__A1 _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07093_ _00614_ _00618_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06605__A2 _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07802__B2 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06044_ _04843_ _04865_ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08358__A2 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05935__I _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09803_ net47 net128 _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07030__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ _00915_ _00855_ _01550_ _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09307__A1 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09734_ _03440_ _03344_ _03349_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06946_ _00371_ _00381_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09858__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09665_ _03276_ _03363_ _03364_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07869__A1 _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06877_ _00396_ _00392_ _00403_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08616_ net111 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08530__A2 _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05828_ _02683_ _02726_ _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09596_ _03270_ _03289_ _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11417__A2 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08547_ _02148_ _02150_ _00674_ net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05759_ net77 _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07097__A2 _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08478_ _02028_ _02030_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07429_ _00758_ _00754_ _00865_ _00741_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10440_ _04176_ _04207_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10371_ _00762_ _04111_ _04133_ net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07546__B _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05845__I _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09010__A3 _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11105__A1 _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06532__A1 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09052__I _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10198__I _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10616__B1 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__A1 _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__B2 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06296__B1 _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10707_ _04424_ _04458_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06835__A2 _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10638_ _04354_ _04385_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09001__B _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07300__I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09785__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10569_ _04317_ _04321_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10395__A2 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11344__A1 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09227__I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07012__A2 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06800_ _00286_ _00327_ _00328_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07780_ _01310_ _01317_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 Operation[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06731_ _00253_ _00260_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09450_ _03093_ _03131_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06662_ _03553_ _05328_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08401_ _01826_ _01942_ _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09381_ _02420_ _01493_ _00968_ _02306_ _03056_ _02546_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_06593_ _00123_ _00124_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08332_ _00780_ _00835_ _00850_ _00774_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08276__A1 _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08263_ _01840_ _01842_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07214_ _00737_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08194_ _00936_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07210__I _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08579__A2 _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07145_ _05665_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07076_ _00556_ _00558_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06027_ _04745_ _04767_ _04865_ _04887_ _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input44_I a_operand[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08200__A1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07978_ _01460_ _01462_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09717_ net126 _02233_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06929_ _00452_ _00456_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_28_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09700__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09648_ _02274_ _01738_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10846__B1 _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06514__A1 _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10310__A2 _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output200_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09579_ _02327_ _02348_ _03176_ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09059__A3 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06278__B1 _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06817__A2 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07490__A2 _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07120__I _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10423_ _03821_ _03925_ _04157_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09767__A1 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10377__A2 _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10354_ _04112_ _04113_ _04114_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_83_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10285_ _03862_ _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11326__A1 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10301__A2 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10656__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06808__A2 _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09758__A1 _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10368__A2 _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07784__A3 _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08981__A2 _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ _02559_ _02571_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11317__A1 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07901_ _01440_ _01448_ _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08881_ _02514_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07832_ _00884_ _01087_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06744__A1 _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07763_ _00815_ _00753_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09502_ _03125_ _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06714_ _05294_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08497__A1 _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07694_ _00819_ _01223_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09433_ net121 net50 _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06645_ net84 net18 _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09364_ _03036_ _03037_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06576_ _05554_ _00106_ _00107_ _00006_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08315_ _01802_ _01897_ _01898_ _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10056__A1 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08464__C _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09295_ _02817_ _01410_ _02962_ _02692_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08246_ net74 net16 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09749__A1 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11005__B1 _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08177_ _01334_ _01050_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07128_ _00463_ _00653_ _00564_ _00562_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07059_ _00416_ _00417_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput160 net160 ALU_Output[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput171 net171 ALU_Output[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput182 net182 ALU_Output[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output150_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput193 net193 ALU_Output[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_43_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10070_ _03742_ _03806_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09516__A4 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08724__A2 _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06735__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10972_ _04618_ _04692_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08488__A1 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10295__A1 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10047__A1 _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09988__A1 _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10598__A2 _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10406_ _03979_ _04169_ _04053_ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11386_ _05225_ _05232_ _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10337_ _04096_ _04066_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10268_ _04018_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10199_ _03833_ _03943_ _03843_ _03946_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__10522__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10286__A1 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06430_ _05609_ _05612_ _05639_ _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05701__A2 _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06361_ _05558_ _05571_ _05572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10589__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08100_ _00775_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09080_ _02659_ _02729_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07454__A2 _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06292_ _05383_ _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08031_ _00795_ _00925_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput40 a_operand[41] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput51 a_operand[51] net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput62 a_operand[61] net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput73 b_operand[13] net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08403__A1 _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput84 b_operand[23] net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput95 b_operand[33] net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08954__A2 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _03504_ _03710_ _03623_ _03624_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _02517_ _02570_ _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08864_ _02402_ _00233_ _00414_ _02381_ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10513__A2 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07815_ _01237_ _01285_ _01321_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_85_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08795_ _02420_ _02292_ _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_38_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07746_ _01279_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07677_ _00901_ _01007_ _01204_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09416_ _03009_ _03012_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06628_ _00086_ _00098_ _00158_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09347_ _03004_ _03018_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06559_ _05408_ _05628_ _03193_ _05477_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ _02864_ _02869_ _02942_ _02941_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__08642__A1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output198_I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08229_ net9 _00766_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11240_ _05058_ _05074_ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09198__A2 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11171_ _04763_ _04990_ _04904_ _04901_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10122_ _03861_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06014__I _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10053_ _03701_ _03719_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09122__A2 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10955_ _04760_ _04764_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10886_ _04512_ _03920_ _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08633__A1 _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05998__A2 _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11369_ _05209_ _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10743__A2 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05930_ _02161_ _02258_ _03813_ _03835_ _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_140_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05861_ _02780_ _02834_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ _01803_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08580_ _01999_ _02186_ _02092_ _02090_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05792_ _02302_ _02335_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_81_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07531_ _01049_ _01050_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07124__A1 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06594__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07462_ _05387_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07675__A2 _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09201_ _02858_ _02859_ _02860_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06413_ _05620_ _05621_ _05622_ _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_50_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07393_ _00915_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09132_ _02362_ _02370_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06344_ _05466_ _05554_ _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09063_ _02592_ _02673_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06275_ _04822_ _02553_ _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05938__I _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10982__A2 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08014_ _01494_ _01486_ _01502_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08927__A2 _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09965_ _02287_ _02326_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08916_ _02540_ _02545_ _02551_ _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09896_ _03613_ _03616_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08847_ _02476_ _02477_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_45_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08778_ net114 _02402_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09104__A2 _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07729_ _01192_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10740_ _04525_ _04529_ _04531_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07666__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08863__A1 _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06874__B1 _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ _04425_ _04451_ _04457_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_13_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06009__I _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__A2 _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05848__I _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11223_ _04996_ _05007_ _05055_ _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09040__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06929__A1 _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10725__A2 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11154_ _04900_ _04905_ _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_122_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10105_ _03842_ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11085_ _04768_ _04774_ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06679__I _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09343__A2 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10036_ _03686_ _03692_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_76_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10489__A1 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10489__B2 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10938_ _04699_ _04711_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07303__I _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10869_ _04587_ _04600_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__A2 _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05758__I _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06093__A1 _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06060_ _05202_ _05234_ _05245_ _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05840__A1 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09582__A2 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__A1 _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09750_ _02977_ _03439_ _03451_ _03458_ net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06962_ _03553_ _02575_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08701_ net119 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05913_ _03651_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09681_ _03296_ _03299_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06893_ _00240_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07345__A1 _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11141__A2 _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08632_ _02238_ _01662_ _01738_ _02240_ _02224_ _02242_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_94_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05844_ _02899_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08563_ _02126_ _02165_ _02167_ _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05775_ _02129_ _02151_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07514_ _04193_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input109_I b_operand[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08494_ _02090_ _02092_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07445_ _05506_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06320__A2 _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07376_ _00890_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09115_ _02719_ _02734_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06327_ _05465_ _05536_ _05537_ _05538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08073__A2 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09270__A1 _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input74_I b_operand[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09046_ _02349_ _02407_ _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06258_ _05411_ _05468_ _05469_ _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09022__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06189_ _05401_ _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08979__I _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07584__A1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09948_ _02387_ _03671_ _03673_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09325__A2 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09879_ _02285_ _02338_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09628__A3 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07639__A2 _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10723_ _04512_ _04309_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06847__B1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06311__A2 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10654_ _04192_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10585_ _04289_ _04363_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09261__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09261__B2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08889__I _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11206_ _05026_ _04171_ _05032_ _05037_ _05038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09564__A2 _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11137_ _04008_ _03932_ _04123_ net44 _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11068_ _04883_ _04886_ _04888_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_49_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10019_ _03747_ _03749_ _03750_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08827__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07230_ _00753_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07161_ _00634_ _00638_ _00685_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06112_ net17 _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10937__A2 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07092_ _00615_ _00617_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07802__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06043_ _05028_ _05060_ _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_114_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09555__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06369__A2 _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11362__A2 _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09802_ net63 net112 _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07994_ _00737_ _00792_ _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09307__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06945_ _00360_ _00471_ _00472_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09733_ _02265_ _02270_ _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06112__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07318__A1 _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11114__A2 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09664_ _03281_ _03333_ _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07869__A2 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06876_ _00403_ _00396_ _00392_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_54_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08467__C _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08615_ _02223_ _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05827_ _02715_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09595_ _02298_ _02355_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06541__A2 _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08546_ _00671_ _02149_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05758_ _01966_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08477_ _01916_ _02029_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09579__B _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09491__A1 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05689_ _01216_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07428_ _01836_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07359_ _00881_ _00875_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09243__A1 _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10928__A2 _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10370_ _00244_ _04122_ _04126_ _02580_ _04132_ _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_109_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09029_ _02670_ _02674_ _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10313__B1 _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10616__A1 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10616__B2 _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10706_ _04424_ _04458_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06296__B2 _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10637_ _04419_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09234__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10568_ _04288_ _04343_ _04345_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09785__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10499_ _04253_ _04270_ _04271_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11344__A2 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06220__A1 _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 a_operand[0] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06730_ _00255_ _00259_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_77_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06867__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06661_ _03465_ _05382_ _00094_ _00191_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_25_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07720__A1 _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08400_ _01950_ _01961_ _01990_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09380_ _02420_ _02964_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06592_ _00052_ _00046_ _00056_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08331_ _01807_ _01916_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06287__A1 _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08262_ _01259_ _01835_ _01841_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06826__A3 _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07213_ _00736_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09225__A1 _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08193_ _00138_ _01679_ _01766_ net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07144_ _00592_ _00669_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07075_ _00453_ _00557_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06026_ _04442_ _04876_ _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input37_I a_operand[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07977_ _01440_ _01448_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09716_ _03417_ _03419_ _03420_ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06928_ _00454_ _00455_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05681__I _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09700__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09647_ _02751_ _03344_ _03345_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10846__B2 _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06859_ _00324_ _00387_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09578_ _03098_ _03270_ _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08529_ _00774_ _01072_ _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08019__A2 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10422_ _04186_ _04187_ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07778__A1 _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10353_ _03825_ _03935_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09519__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10284_ _03860_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11326__A2 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06202__A1 _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06269__A1 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11262__A1 _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10065__A2 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07311__I _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09207__A1 _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11014__A1 _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09758__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07769__A1 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05766__I _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06441__A1 _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07900_ _01443_ _01447_ _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08880_ net50 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07831_ _01310_ _01317_ _01372_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10621__B _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05715__B _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06597__I _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07762_ _01049_ _00806_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09143__B1 _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09501_ _03122_ _03123_ _03126_ _03029_ _03027_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_37_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06713_ _00210_ _00237_ _00222_ _00238_ _00242_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07693_ net91 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08497__A2 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09432_ _03026_ _03031_ _03035_ _03111_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_25_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06644_ _00007_ _00173_ _00174_ _00109_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_24_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09363_ _03031_ _03035_ _03026_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06575_ _00003_ _00007_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08249__A2 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08314_ _01805_ _01818_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10056__A2 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09997__A2 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09294_ _02961_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08245_ _00778_ _01161_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11005__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08176_ _01647_ _01746_ _01747_ _01545_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_21_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07127_ _02280_ _03411_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05676__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07058_ _00584_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput150 net150 ALU_Output[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_133_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput161 net161 ALU_Output[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput172 net172 ALU_Output[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06009_ _04691_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xoutput183 net183 ALU_Output[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_102_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput194 net194 ALU_Output[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output143_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06300__I _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10971_ _04780_ _04781_ _04782_ _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08488__A2 _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10295__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09437__A1 _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10047__A2 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07999__A1 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08948__B1 _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10405_ _03975_ _03978_ _03942_ _03969_ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_109_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11385_ _05227_ _05229_ _05231_ _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08412__A2 _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10336_ _03827_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ _04018_ _04020_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10198_ _03945_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07306__I _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10286__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09140__A3 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09428__A1 _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11235__A1 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06360_ _05564_ _05570_ _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10038__A2 _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06291_ _05502_ _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08030_ _00926_ _01503_ _01504_ _00795_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06662__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput30 a_operand[32] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput41 a_operand[42] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput52 a_operand[52] net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput63 a_operand[62] net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_116_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput74 b_operand[14] net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput85 b_operand[24] net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09600__A1 _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput96 b_operand[34] net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_66_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06414__A1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ _02300_ _03006_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08932_ _02562_ _02566_ _02569_ _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08863_ _02483_ _02254_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07814_ _01353_ _01327_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08794_ _02287_ _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07745_ _01209_ _01245_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07676_ _01007_ _01203_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09415_ _03020_ _03091_ _03092_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09419__A1 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06627_ _00087_ _00097_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08890__A2 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11226__A1 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09346_ _03013_ _03017_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06558_ _00077_ _00088_ _00089_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09277_ _02939_ _02941_ _02942_ _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06489_ _05381_ _00018_ _00021_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_32_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08642__A2 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06653__A1 _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08228_ _01725_ _01732_ _01804_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _00805_ _01157_ _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06405__A1 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11170_ _04774_ _04997_ _04998_ _04331_ _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_107_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10121_ net42 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08158__A1 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10052_ _03703_ _03718_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07905__A1 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__B1 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06030__I _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09122__A3 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10954_ _04761_ _04762_ _04763_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_16_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08330__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10885_ _03886_ _03912_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_16_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05695__A2 _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08633__A2 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07796__I _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06644__A1 _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11368_ _05211_ _05214_ _00674_ net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10319_ _04074_ _04077_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11299_ _05138_ _05107_ _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07464__C _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09897__A1 _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05860_ _02780_ _02834_ _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10900__B1 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05791_ _02324_ _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09649__A1 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10259__A2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07530_ _00877_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07480__B _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07124__A2 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08295__C _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07461_ _01640_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06412_ _02543_ _05126_ _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09200_ _02220_ _02309_ _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07392_ _00914_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09131_ _02779_ _02781_ _02784_ _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06343_ _02478_ _05413_ _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09062_ _02649_ _02708_ _02709_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10431__A2 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06274_ _05466_ _05470_ _05485_ _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08013_ _01511_ _01570_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10719__B1 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06115__I _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09964_ _02296_ _02314_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05954__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09337__B1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08915_ _02382_ _02391_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09895_ _03614_ _03615_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_85_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08846_ net48 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08560__A1 _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08777_ _02387_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05989_ _04086_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07728_ _01261_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07115__A2 _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07659_ _00045_ _01186_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06874__A1 _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10670__A2 _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10670_ _04452_ _04454_ _04456_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__06874__B2 _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09329_ _02936_ _02946_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06626__A1 _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11222_ _04980_ _04994_ _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09040__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11153_ _04900_ _04905_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07565__B _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05864__I _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ _03841_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11084_ _04894_ _04900_ _04905_ _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09879__A1 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10035_ _03764_ _03767_ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10489__A2 _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07106__A2 _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10937_ _04096_ _03854_ _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07657__A3 _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10661__A2 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10868_ _04597_ _04610_ _04670_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09803__A1 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10799_ _04529_ _04531_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10964__A3 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06093__A2 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08790__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06961_ _00269_ _00480_ _00369_ _00366_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08700_ _02311_ _02316_ _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05912_ _03640_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09680_ _03296_ _03299_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06892_ _00416_ _00417_ _00238_ _00419_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08631_ _01825_ _02241_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05843_ _02889_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08562_ _00931_ _01072_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05774_ _02140_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ _00881_ _00211_ _00212_ _00967_ _01033_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10101__A1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08493_ _02087_ _02091_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07648__A3 _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07444_ _00847_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07375_ _00887_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09114_ _02713_ _02714_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06326_ _05462_ _05492_ _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_109_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09270__A2 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06257_ _05467_ _05417_ _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06084__A2 _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09045_ _01192_ _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input67_I a_operand[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06188_ _05346_ _05371_ _05401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09022__A2 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07033__A1 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09156__I _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05684__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07584__A2 _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09947_ _02479_ _02256_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09878_ _02295_ _02323_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08829_ _02282_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10340__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08297__B1 _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10722_ net103 _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10643__A2 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10653_ _04234_ _03937_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10584_ _03877_ _04231_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09261__A2 _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11205_ _00959_ _05033_ _05034_ _05036_ _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11136_ _04880_ _04960_ _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11067_ _03872_ _04439_ _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08524__A1 _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10018_ _03586_ _03747_ _03749_ _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10882__A2 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08827__A2 _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07160_ _00631_ _00684_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09252__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06111_ _05279_ _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07091_ _00612_ _00616_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06042_ _05039_ _05049_ _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ _03417_ _03513_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06369__A3 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07993_ _01535_ _01548_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_86_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09732_ _03360_ _03435_ _03438_ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_39_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06944_ _00365_ _00370_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09663_ _03281_ _03333_ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06875_ _02096_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input121_I b_operand[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08614_ _02222_ _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05826_ _02704_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09594_ _03287_ _02370_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08545_ _02065_ _02147_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05757_ _01390_ _01944_ _01955_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06829__A1 _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ _02024_ _02071_ _02072_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05688_ _01205_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09491__A2 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ _05497_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05679__I _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07358_ _00872_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06309_ _05434_ _05517_ _05520_ _05449_ _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07289_ _00811_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09028_ _02591_ _02673_ _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_output173_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06303__I _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10561__A1 _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10561__B2 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06517__B1 _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10313__A1 _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10616__A2 _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _04487_ _04491_ _04492_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06296__A2 _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07493__A1 _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10636_ _04356_ _04417_ _04418_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10567_ _04285_ _04322_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_10_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10498_ _01477_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07309__I _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11119_ _04878_ _04891_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 a_operand[10] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10855__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06660_ _03455_ _05408_ _05412_ _03367_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06591_ _00052_ _00046_ _00056_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_33_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ net9 _00834_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08261_ _00906_ _00892_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07484__A1 _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07212_ net5 _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08192_ _01680_ _01682_ _01691_ _01765_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09225__A2 _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07236__A1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07143_ _00665_ _00668_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08984__A1 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07074_ _00552_ _00598_ _00599_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10791__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06025_ _04843_ _04854_ _04420_ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07219__I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10543__A1 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07976_ _01449_ _01465_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09434__I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09715_ _03326_ _03416_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_74_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06927_ _02172_ _02824_ _02965_ net26 _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09646_ _03239_ _03249_ _03230_ _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_83_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09700__A3 _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06858_ _00326_ _00386_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10846__A2 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07711__A2 _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05809_ net20 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09577_ net56 _02344_ _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06789_ _00247_ _00248_ _00306_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08528_ _01927_ _02130_ _02037_ _02035_ _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_70_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07475__A1 _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08459_ _01853_ _01969_ _01970_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_51_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08019__A3 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _03822_ _03915_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08975__A1 _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10352_ _03959_ _03842_ _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10283_ _03852_ _03855_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06202__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05872__I _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05961__A1 _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07702__A2 _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06269__A2 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10619_ _04400_ _01651_ _00126_ _04028_ _04401_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07769__A2 _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10525__A1 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07830_ _01313_ _01316_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07761_ _01289_ _01293_ _01296_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09500_ _03173_ _03185_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_49_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06712_ _05380_ _00239_ _00241_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07692_ _00870_ _00833_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09431_ _03032_ _03034_ _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06643_ _00106_ _00110_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09362_ _03026_ _03031_ _03035_ _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06574_ _02412_ _05353_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09446__A2 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08313_ _01805_ _01818_ _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_32_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09293_ _02296_ _02300_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08244_ _01048_ _00933_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11005__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08175_ _00810_ _00889_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10213__B1 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08957__A1 _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ _00649_ _00651_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10764__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10764__B2 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06432__A2 _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07057_ _05387_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput140 net140 ALU_Output[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput151 net151 ALU_Output[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput162 net162 ALU_Output[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06008_ _03988_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput173 net173 ALU_Output[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput184 net184 ALU_Output[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10516__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput195 net195 ALU_Output[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06196__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05692__I _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07959_ _01438_ _01475_ _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output136_I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10103__I _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ _04707_ _04710_ _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06499__A2 _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07696__A1 _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09629_ _03201_ _03326_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09437__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07412__I _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07448__A1 _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06120__A1 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06120__B2 _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08948__A1 _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _04052_ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08948__B2 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11384_ _05188_ _05228_ _05230_ _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_137_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10755__A1 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10335_ _04076_ _04094_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10266_ _04019_ _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10197_ _03814_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05934__A1 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09140__A4 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09428__A2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07322__I _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11235__A2 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06290_ _04075_ _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 a_operand[23] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput31 a_operand[33] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput42 a_operand[43] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05777__I _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput53 a_operand[53] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08939__A1 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput64 a_operand[63] net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput75 b_operand[15] net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput86 b_operand[25] net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_143_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09600__A2 _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput97 b_operand[35] net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09980_ _03704_ _03708_ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08931_ _02488_ _02518_ _02568_ _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08167__A2 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08862_ _05375_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07914__A2 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07813_ _01284_ _01322_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08793_ _02307_ _02317_ _02418_ _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07744_ _01273_ _01276_ _01976_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07675_ _01143_ _01146_ _01202_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09414_ _03021_ _03036_ _03037_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06626_ _04107_ _02183_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06350__A1 _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09419__A2 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07232__I _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09345_ _02746_ _03015_ _03016_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_52_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11226__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06557_ _02357_ _02943_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input97_I b_operand[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09276_ _02229_ _02301_ _02315_ _02251_ _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06488_ _03433_ _03258_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ _01728_ _01731_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06653__A2 _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08158_ net130 _00892_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10737__A1 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07109_ _03694_ _02596_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07602__A1 _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06405__A2 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08089_ _01635_ _01653_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10120_ _03859_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08158__A2 _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10051_ _03780_ _03782_ _03785_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_76_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11162__A1 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09107__A1 _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09107__B2 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07669__A1 _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ net106 _03956_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09122__A4 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08330__A2 _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10884_ _04513_ _04686_ _04687_ _04623_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__06341__A1 _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08094__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10976__A1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07841__A1 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06644__A2 _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10728__A1 _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09594__A1 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11367_ _00671_ _05212_ _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10318_ _03828_ _03844_ _04076_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08701__I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11298_ _05089_ _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08149__A2 _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10249_ _03860_ _03863_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11153__A1 _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09897__A2 _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10900__A1 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05790_ _02313_ _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09649__A2 _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06580__A1 _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08321__A2 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07460_ _00979_ _00980_ _00981_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08148__I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06411_ _03564_ _01998_ _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07391_ _00913_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09130_ _02671_ _02783_ _02333_ _02234_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__08085__A1 _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06342_ _02596_ _01585_ _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10967__A1 _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10627__B _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09061_ _02652_ _02676_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06273_ _05484_ _05485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07832__A1 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06635__A2 _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10431__A3 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08012_ _01514_ _01569_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10719__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10719__B2 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10195__A2 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08611__I _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09963_ _03523_ _03676_ _03587_ _03588_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08914_ _02520_ _02523_ _02534_ _02550_ net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09894_ _02432_ _02356_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11144__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ _02248_ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08560__A2 _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08776_ _02231_ _02253_ _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06571__A1 _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05988_ _04054_ _04139_ _04225_ _04464_ net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input12_I a_operand[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07727_ _01259_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11193__B _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10655__B1 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07658_ _01117_ _01128_ _01144_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06609_ _00139_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07589_ _01081_ _01110_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09328_ _02919_ _02933_ _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08076__A1 _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10958__A1 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ _02920_ _02922_ _02923_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11221_ _04979_ _05009_ _05053_ _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11152_ _04955_ _04958_ _04978_ _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__11368__B _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10103_ _03840_ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11083_ _04901_ _04904_ _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11135__A1 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09879__A2 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08000__A1 _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10034_ _02961_ _03765_ _03766_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_49_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08551__A2 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06562__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05880__I _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10498__I _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10936_ _04677_ _04716_ _04743_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06314__A1 _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10867_ _04598_ _04609_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08067__A1 _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10798_ _04529_ _04531_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10949__A1 _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08606__A3 _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09803__A2 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07600__I _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11419_ _05259_ _05263_ _05269_ _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_125_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09031__A3 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06960_ _00279_ _00486_ _00487_ _05514_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I Operation[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05911_ net87 _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06891_ _00418_ _00416_ _00417_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08630_ _02240_ _01890_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05842_ net14 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07491__B _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06886__I _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08561_ _02036_ _02165_ _02134_ _02132_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05773_ net90 _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07512_ _01346_ _00841_ _01032_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__10201__I _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08492_ net74 _00828_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10101__A2 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07443_ _04626_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10652__A3 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07374_ _00891_ _00896_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09113_ _02740_ _02742_ _02764_ _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06325_ _05462_ _05492_ _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09044_ _04485_ _02689_ _02690_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06256_ _05467_ _05417_ _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06187_ _05394_ _05398_ _05292_ _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08230__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07033__A2 _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09946_ _02260_ _02386_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09877_ _03423_ _03584_ _03595_ _03522_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_85_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08828_ _02278_ _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__I _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08759_ _02245_ _02239_ _02252_ _02381_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09494__B1 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08297__B2 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10721_ _03886_ _04307_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06847__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10652_ _04434_ _04435_ _04436_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10583_ _03890_ _03816_ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09549__A1 _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__B2 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11204_ _04842_ _05026_ _04593_ _05035_ _05036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_122_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11135_ net44 _04183_ _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08772__A2 _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11108__A1 _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06783__A1 _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11066_ _04701_ _04306_ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08524__A2 _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ _02264_ _02581_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10331__A2 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07732__B1 _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10619__B1 _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08288__A1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06838__A2 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ _04725_ _04726_ _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07330__I _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07799__B1 _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06110_ _05324_ _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07090_ net92 _02748_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06041_ net76 _02769_ _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10691__I _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06471__B1 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11347__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05785__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09800_ _03417_ _03419_ _03420_ _03426_ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07992_ _01536_ _01547_ _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09731_ _03436_ _03437_ _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06943_ _00365_ _00370_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08515__A2 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09712__A1 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _03268_ _03274_ _03361_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06874_ _05446_ _00316_ _00390_ _05496_ _00402_ net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_28_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08613_ _02221_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05825_ _02694_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09593_ _02289_ _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input114_I b_operand[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08544_ _02065_ _02147_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08279__A1 _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05756_ _01433_ _01444_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10086__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08475_ _02070_ _02040_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05687_ _01162_ _01195_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07426_ _00769_ _00948_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ _00821_ _00826_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08780__B _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06308_ _05519_ _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07288_ _00810_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10815__B _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09027_ _02671_ _02347_ _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06239_ _05393_ _05396_ _05450_ _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07006__A2 _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output166_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09951__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06765__A1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10561__A2 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09929_ _02444_ _02443_ _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08506__A2 _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06517__A1 _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08911__C1 _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10704_ _04487_ _04491_ _03254_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07493__A2 _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07150__I _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10635_ _04351_ _04315_ _04359_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_127_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10566_ _04285_ _04322_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08442__A1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10497_ _03918_ _03980_ _04108_ _04268_ _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11118_ _04878_ _04891_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11049_ _04096_ _04019_ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 a_operand[11] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10304__A2 _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07325__I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__A1 _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06590_ _00062_ _00121_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05731__A2 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08260_ _01552_ _01829_ _01839_ _01717_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07211_ _00675_ _00732_ _00733_ _00735_ net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08191_ _00992_ _01764_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07142_ _00508_ _00666_ _00667_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06444__B1 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08984__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07073_ _00597_ _00567_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10791__A2 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06024_ _04420_ _04843_ _04854_ _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_126_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09933__A1 _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06211__A3 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07975_ _01521_ _01528_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09714_ _02275_ _02563_ _03418_ _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06926_ _00347_ _00453_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09161__A2 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09645_ _03239_ _03230_ _02464_ _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06857_ _00336_ _00385_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05808_ _02467_ _02510_ _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09576_ _03173_ _03185_ _03267_ _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06788_ _00149_ _00204_ _00309_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08527_ _00790_ _00890_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05739_ _01760_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08458_ _01776_ _02054_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07475__A2 _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07409_ _00931_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08389_ _01906_ _01978_ _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10420_ _04156_ _04181_ _04185_ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10351_ _03952_ _03815_ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08975__A2 _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08015__B _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10782__A2 _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10282_ _04037_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09924__A1 _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05961__A2 _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10298__A1 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07702__A3 _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06910__A1 _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08663__A1 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08704__I _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10618_ _04335_ _04279_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10222__A1 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10549_ _04030_ _04255_ _04259_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_116_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09915__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10525__A2 _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07760_ _01294_ _01295_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06711_ _03824_ _00240_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07691_ _00885_ _00765_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09430_ _03096_ _03109_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06642_ net86 _05213_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06901__A1 _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _03032_ _03034_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06573_ _00101_ _00104_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08103__B1 _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08312_ _01894_ _01895_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09292_ _02958_ _02959_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_61_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08243_ _01714_ _01720_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08174_ _00896_ _01648_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10213__A1 _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07125_ _00557_ _00650_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10213__B2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08957__A2 _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10764__A2 _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07056_ _00577_ _00582_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput141 net141 ALU_Output[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput152 net152 ALU_Output[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06007_ _03041_ _03052_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09906__A1 _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput163 net163 ALU_Output[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput174 net174 ALU_Output[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input42_I a_operand[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10516__A2 _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput185 net185 ALU_Output[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput196 net196 ALU_Output[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07958_ _01508_ _01510_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06909_ _00345_ _00357_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07889_ _01393_ _01397_ _01435_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09628_ _02227_ net62 _02432_ _02250_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09559_ _02431_ _02438_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10452__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06120__A2 _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10403_ _04031_ _03973_ _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08948__A2 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11383_ _04020_ _03975_ _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10334_ _03820_ _03951_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10265_ net45 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10196_ _03822_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05934__A2 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07439__A2 _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08636__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10443__A1 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 a_operand[14] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput21 a_operand[24] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput32 a_operand[34] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 a_operand[44] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput54 a_operand[54] net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput65 a_operand[6] net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput76 b_operand[16] net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10746__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput87 b_operand[26] net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput98 b_operand[36] net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07611__A2 _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08930_ _02567_ _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06889__I _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05793__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08861_ _02475_ _00421_ _02482_ _04604_ _02493_ _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06178__A2 _05391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08102__C _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07914__A3 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07812_ _01347_ _01351_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08792_ _02330_ _02415_ _02416_ _02417_ _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07743_ _01273_ _01276_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07127__A1 _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07674_ _00898_ _00899_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06625_ _00081_ _00115_ _00155_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09413_ _03036_ _03037_ _03021_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06350__A2 _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09344_ _02326_ _02392_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06556_ net23 net77 _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10434__A1 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09275_ _02507_ _02940_ _02937_ _02938_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_138_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06487_ _05568_ _00018_ _00019_ _05627_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08226_ _01745_ _01800_ _01801_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08157_ _01550_ _01715_ _01726_ _01622_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07108_ _00632_ _00633_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08088_ _01638_ _01652_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07602__A2 _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07039_ _00561_ _00565_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ _03783_ _03784_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11162__A2 _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10114__I _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10370__B1 _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__A2 _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10952_ net105 net33 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07669__A2 _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10883_ _04620_ _04624_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06341__A2 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09291__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10976__A2 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07841__A2 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09043__A1 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09594__A2 _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11366_ _05131_ _05210_ _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10317_ _03961_ _03816_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11297_ _05106_ _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10248_ _03875_ _03986_ _03997_ _04000_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10179_ _03924_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07109__A1 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06580__A2 _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06410_ _05560_ _05302_ _05620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08609__A1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07390_ net70 _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10416__A1 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06341_ _01108_ _02500_ _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05788__I _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09060_ _02652_ _02676_ _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06272_ _05475_ _05483_ _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07832__A2 _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10431__A4 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08011_ _01516_ _01519_ _01568_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_135_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10719__A2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09962_ _03687_ _03688_ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07508__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08913_ _02495_ _02538_ _02549_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09893_ _02279_ _03387_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11144__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08844_ _02252_ _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08775_ _02382_ _02391_ _02397_ _02398_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_05987_ _01141_ _04269_ _04355_ _04453_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_27_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06571__A2 _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07726_ net66 net130 _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07243__I _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10655__B2 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07657_ _01144_ _01117_ _01128_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_41_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06608_ _02205_ _02247_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07588_ _01083_ _01109_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06539_ _00001_ _00026_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09327_ _02992_ _02996_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08076__A2 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09273__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05698__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11080__A1 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09258_ _02351_ _02359_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output196_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08209_ _01710_ _01756_ _01783_ _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09189_ _02843_ _02847_ _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09025__A1 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10109__I _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11220_ _04985_ _05008_ _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08802__I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11383__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11151_ _04965_ _04977_ _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10591__B1 _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10102_ net95 _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11082_ _04902_ _04903_ _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10033_ _02259_ _02393_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08000__A2 _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10894__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10935_ _04681_ _04715_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07511__A1 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10866_ _04096_ _04008_ _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09264__A1 _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08067__A2 _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10797_ _04507_ _04515_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09016__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11418_ _05264_ _05266_ _05268_ _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07578__A1 _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11349_ _03854_ _03924_ _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06232__I _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11126__A2 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05910_ net23 _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06890_ _01944_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05841_ _02867_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07750__A1 _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08560_ _00781_ _00899_ _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05772_ _02118_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07511_ _01944_ _01031_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08491_ _00777_ _01102_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09699__B _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07998__I _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07442_ _00955_ _00963_ _00964_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07373_ _00893_ _00895_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06069__A1 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06324_ _05456_ _05457_ _05494_ _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09112_ _02706_ _02739_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09043_ _02627_ _02637_ _02688_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_06255_ _05301_ _05414_ _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06186_ _05394_ _05398_ _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09022__A4 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08230__A2 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09945_ _03668_ _03669_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09876_ _03521_ _03523_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08827_ _02263_ _02268_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08758_ _02380_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07709_ _00842_ _01159_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08297__A2 _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09494__A1 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08689_ _02297_ _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09494__B2 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10720_ _04361_ _04508_ _04509_ _04426_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10651_ _03893_ _03950_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10582_ _04191_ _03879_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06317__I _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07857__B _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09549__A2 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11203_ _05202_ _03847_ _05026_ _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07148__I _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11134_ net45 _04295_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11065_ _04709_ _04883_ _04884_ _04795_ _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_62_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10016_ _03238_ _02621_ _03678_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_76_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07732__A1 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10302__I _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10619__A1 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10619__B2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10918_ _04641_ _04723_ _04722_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08707__I _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09237__A1 _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10849_ _04930_ _04565_ _04639_ _04650_ net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__11044__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09788__A2 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07799__A1 _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07799__B2 _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06040_ _01108_ _02976_ _01564_ _02020_ _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__11289__B _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06471__B2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11347__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07058__I _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ _01539_ _01543_ _01546_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_68_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07971__A1 _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09730_ _03261_ _03337_ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06942_ _00448_ _00451_ _00469_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__06897__I _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05982__B1 _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09661_ _02459_ _02540_ _03275_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09712__A2 _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06873_ _00391_ _00393_ _00401_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08612_ _02220_ _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05824_ net82 _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09592_ _03194_ _03198_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08543_ _02143_ _02146_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05755_ _01401_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input107_I b_operand[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09222__B _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08474_ _02070_ _02040_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05686_ _01173_ _01184_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07425_ _00747_ _00945_ _00947_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07356_ _00876_ _00878_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06307_ _05518_ _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07287_ _00809_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input72_I b_operand[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06462__A1 _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09026_ _02219_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06238_ _03498_ _03509_ _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06169_ _01618_ _01694_ _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10010__A2 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09951__A2 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output159_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09928_ _00671_ _03652_ _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09164__B1 _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09703__A2 _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10849__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09859_ _03519_ _03524_ _03576_ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06517__A2 _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08911__B1 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10313__A3 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10122__I _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08911__C2 _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07431__I _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10703_ _03875_ _03986_ _04055_ _04490_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09219__A1 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10634_ _04351_ _04315_ _04359_ _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06047__I _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10565_ _04284_ _04340_ _04341_ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05886__I _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10496_ _04265_ _04051_ _04267_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06205__A1 _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11117_ _04938_ _04939_ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09093__I _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11048_ _04861_ _04866_ _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 a_operand[12] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__A2 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08130__A1 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06141__B1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07210_ _00734_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08190_ _01693_ _01763_ _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06692__A1 _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07141_ _00512_ _00571_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09630__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05796__I _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06444__A1 _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ _00597_ _00567_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06023_ _04800_ _04811_ _04832_ _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06995__A2 _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10207__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09933__A2 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06747__A2 _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07974_ _01523_ _01527_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09713_ _02793_ _02266_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06925_ net26 _02824_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09644_ _00244_ _03342_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06856_ _00340_ _00384_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05807_ _02500_ _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09575_ _03174_ _03184_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06787_ _03922_ _00315_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08526_ _02125_ _02127_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05738_ _01749_ _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07251__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08121__A1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08457_ _01887_ _01969_ _02052_ _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07408_ net10 _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06683__A1 _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08388_ _01965_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07339_ _00856_ _00857_ _00861_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06435__A1 _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10350_ _03967_ _04110_ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06986__A2 _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09009_ _02516_ _02567_ _02597_ _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__10117__I _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10281_ _03972_ _04030_ _04036_ _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09924__A2 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08810__I _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09688__A1 _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10298__A2 _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11247__A1 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08663__A2 _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06674__A1 _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10617_ _03874_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09612__A1 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10222__A2 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10548_ _04281_ _04284_ _04324_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_6_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10479_ _04188_ _04205_ _04249_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08720__I _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06710_ _01716_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07690_ _01219_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08351__A1 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06641_ _00102_ _00170_ _00171_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_64_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _03027_ _03029_ _03033_ _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06572_ _00103_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08103__A1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08311_ _01795_ _01849_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09291_ _02891_ _02884_ _02461_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08242_ _01721_ _01733_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08173_ _01742_ _01744_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08406__A2 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09603__A1 _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06417__A1 _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11410__A1 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07124_ _02053_ _02845_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06968__A2 _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07090__A1 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07055_ _00317_ _00580_ _00581_ _00579_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput142 net142 ALU_Output[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06006_ _01596_ _04269_ _04582_ _04604_ _04658_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_82_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput153 net153 ALU_Output[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput164 net164 ALU_Output[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput175 net175 ALU_Output[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07917__A1 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10381__B _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput186 net186 ALU_Output[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput197 net197 Exception[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_43_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input35_I a_operand[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07957_ _01480_ _01482_ _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06908_ _00345_ _00357_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07888_ _01307_ _01395_ _01394_ _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09627_ _03323_ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06839_ net88 _05213_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09558_ _02464_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08509_ _00919_ _00815_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09489_ _03025_ _03116_ _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08645__A2 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06656__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08805__I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10452__A2 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06408__A1 _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10402_ _04136_ _04138_ _04148_ _04166_ net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__11401__A1 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11382_ _05101_ _05228_ _05196_ _05194_ _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10755__A3 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10333_ _03254_ _04092_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10264_ _04017_ _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10195_ _03936_ _03941_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08581__A1 _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06895__A1 _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10979__B1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08636__A2 _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06647__A1 _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput11 a_operand[15] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput22 a_operand[25] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput33 a_operand[35] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput44 a_operand[45] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput55 a_operand[55] net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput66 a_operand[7] net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09061__A2 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput77 b_operand[17] net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput88 b_operand[27] net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput99 b_operand[37] net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09546__I _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08021__B1 _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08860_ _00951_ _02491_ _02492_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_112_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07811_ _01137_ _01349_ _01350_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08791_ _02311_ _02316_ _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07742_ _00818_ _00945_ _01274_ _01275_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_38_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07127__A2 _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07673_ _01200_ _00902_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09412_ _03083_ _03089_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06624_ _00010_ _00025_ _00114_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09343_ _03014_ _02366_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06555_ _00005_ _00008_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09824__A1 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06638__A1 _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09274_ _02299_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06486_ _05360_ _03193_ _05223_ _05477_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08225_ _01748_ _01752_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08156_ _01048_ _00785_ _00792_ _01161_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06145__I _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07063__A1 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07107_ _00532_ _00535_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08087_ _01639_ _01650_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07038_ _00562_ _00564_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output141_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08989_ _02631_ _02447_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10370__A1 _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10370__B2 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08315__A1 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10951_ net107 _03809_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10130__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10882_ _03865_ _04307_ _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09815__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11365_ _05131_ _05210_ _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05894__I _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10316_ _03971_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06801__A1 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11296_ _05133_ _05134_ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10247_ _03998_ _03994_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10178_ _03923_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07109__A2 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09806__A1 _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06340_ _05544_ _05547_ _05550_ _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06271_ _05479_ _05482_ _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08010_ _01529_ _01567_ _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09961_ _03598_ _03600_ _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08912_ _02541_ _02544_ _02548_ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09892_ _02462_ _02392_ _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08843_ _02246_ _02254_ _02473_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07899__A3 _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08774_ _02384_ _02389_ _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05986_ _04388_ _04399_ _04431_ _04442_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07725_ _01256_ _00983_ _01257_ _01199_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06859__A1 _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10655__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ _01181_ _01182_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06607_ _00137_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07587_ _01093_ _01107_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05979__I _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09326_ _02993_ _02995_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06538_ _00028_ _00066_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_139_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09273__A2 _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11080__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ _02452_ _02372_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06469_ _01086_ _03640_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08208_ _01712_ _01755_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09387__S _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _02723_ _02844_ _02846_ _02786_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09025__A2 _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output189_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07036__A1 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08139_ _01641_ _01704_ _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11150_ _04975_ _04976_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10591__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10591__B2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10101_ _03833_ _03832_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10125__I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11081_ net106 _03937_ _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10032_ _02287_ _02315_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06011__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10894__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10646__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10934_ _04671_ _04675_ _04741_ _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07511__A2 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10865_ _04665_ _04666_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05889__I _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10796_ _04518_ _04533_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09264__A2 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09016__A2 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11417_ _03992_ _03880_ _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11348_ _04971_ _05192_ _05102_ _05100_ _05193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_4_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11279_ _05112_ _05117_ _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_140_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08527__A1 _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05840_ _02791_ _02856_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10885__A2 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05771_ _02107_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07510_ _01030_ _00833_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08490_ _01824_ _02087_ _02088_ _01997_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_62_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07441_ _01412_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05799__I _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07372_ _00894_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09111_ _02451_ _02762_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06323_ _05461_ _05493_ _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09042_ _02627_ _02688_ _02636_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06254_ _05300_ _02586_ _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08903__I _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09000__S _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07018__A1 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06185_ _05396_ _05397_ _04702_ _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09944_ _03591_ _03603_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06241__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09875_ _03593_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10325__A1 _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ _02404_ _02449_ _02451_ _02454_ _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_85_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07254__I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08757_ _02235_ _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05752__A1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05969_ _04258_ _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07708_ _01155_ _01167_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ _02297_ _02303_ _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09494__A2 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07639_ _00737_ _00889_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10650_ _03882_ _03840_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09246__A2 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09309_ _02881_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11053__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10581_ _04352_ _04356_ _04359_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_108_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11202_ _03848_ _01418_ _05507_ _04817_ _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11133_ _04910_ _04915_ _04957_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11064_ _04793_ _04796_ _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10015_ _03662_ _03744_ _03745_ _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07732__A2 _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05743__A1 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10619__A2 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09485__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10917_ _04722_ _04641_ _04723_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_71_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06508__I _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10848_ _04040_ _01251_ _04642_ _01255_ _04649_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_20_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11044__A2 _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10779_ _04535_ _04540_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_9_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07799__A2 _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08996__A1 _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08723__I _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06471__A2 _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07990_ _01541_ _01544_ _01545_ _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_87_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06941_ _00457_ _00468_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05982__A1 _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09660_ _03222_ _03223_ _03357_ _03359_ _03340_ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_67_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10858__A2 _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06872_ _00231_ _05180_ _00399_ _00400_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08611_ _02219_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05823_ _02672_ _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09591_ _03282_ _03284_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08542_ _01975_ _02144_ _02145_ _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05754_ _01141_ _01249_ _01509_ _01923_ net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08473_ _02027_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05685_ net2 _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07424_ _00742_ _00758_ _00946_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09228__A2 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07355_ _00871_ _00877_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08987__A1 _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06306_ _01466_ _01673_ _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07286_ net66 _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10794__A1 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09025_ _02393_ _02387_ _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06237_ _05448_ _03542_ _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07249__I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input65_I a_operand[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06168_ _05381_ _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06099_ _03095_ _05147_ _05314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09464__I _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09927_ _03648_ _03649_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09164__A1 _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09164__B2 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09858_ _03575_ _03518_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08911__A1 _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08911__B2 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08809_ _02436_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09789_ _03298_ _03500_ _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09413__B _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _04134_ _04479_ _04489_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10633_ _04350_ _04414_ _04415_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_41_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08978__A1 _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10564_ _04281_ _04324_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07650__A1 _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10495_ _03974_ _03979_ _04169_ _04266_ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_142_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06063__I _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11116_ _04869_ _04921_ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11047_ _04863_ _04864_ _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 a_operand[13] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_49_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08718__I _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09458__A2 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07469__A1 _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08969__A1 _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07140_ _00512_ _00571_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09630__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07071_ _00555_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06444__A2 _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06022_ _04800_ _04811_ _04832_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10528__A1 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08197__A2 _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09394__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06701__I _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07973_ _01454_ _01524_ _01526_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05955__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09712_ _03326_ _03416_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06924_ net28 _02020_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09643_ _03257_ _03341_ _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06855_ _00358_ _00383_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05806_ _02489_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09574_ _02281_ _02384_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08628__I _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06786_ _03845_ _04951_ _00314_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08525_ _02029_ _02126_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05737_ _01281_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10059__A3 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08121__A2 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08456_ _01889_ _01891_ _01968_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07407_ _00779_ _00788_ _00927_ _00929_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08387_ _01908_ _01964_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07880__A1 _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06592__B _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07338_ _00859_ _00860_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_13_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09621__A2 _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07269_ net71 _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09008_ _02594_ _02651_ _02604_ _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output171_I net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10280_ _04031_ _04033_ _04035_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09385__A1 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11192__A1 _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07935__A2 _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09137__A1 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10133__I _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09688__A2 _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11247__A2 _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09860__A2 _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10470__A3 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05897__I _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10616_ _03880_ _00988_ _04395_ _00989_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10547_ _04285_ _04288_ _04322_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07623__A1 _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10478_ _04186_ _04187_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_6_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09376__A1 _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05937__A1 _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10930__A1 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06640_ _01108_ _02237_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06362__A1 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07352__I _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06571_ _00002_ _00102_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_80_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08310_ _01799_ _01848_ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09300__A1 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08103__A2 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09300__B2 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09290_ _02891_ _02957_ _02884_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_61_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06114__A1 _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08241_ _01802_ _01805_ _01818_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_123_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07862__A1 _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06665__A2 _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08172_ _01706_ _01743_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07123_ net28 _02845_ _04539_ _02053_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11410__A2 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07054_ _00389_ _00502_ _00503_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__07090__A2 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06005_ _04301_ _04626_ _04648_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput143 net143 ALU_Output[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput154 net154 ALU_Output[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput165 net165 ALU_Output[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10381__C _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput176 net176 ALU_Output[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput187 net187 ALU_Output[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_141_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput198 net198 Exception[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09119__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10921__A1 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__B2 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07956_ _01434_ _01478_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input28_I a_operand[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06907_ _00433_ _00434_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07887_ _01362_ _01431_ _01432_ _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10685__B1 _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09626_ _02508_ _02462_ _02433_ _02251_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06838_ _02216_ _02889_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07550__B1 _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11229__A2 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09557_ _02977_ _03225_ _03242_ _03247_ net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_43_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06769_ _00295_ _00297_ _00298_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_71_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ _02106_ _02108_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09488_ _03100_ _03108_ _03172_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ _01815_ _02033_ _01928_ _01926_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06656__A2 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07211__B _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06606__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10401_ _02152_ _04165_ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11381_ _04008_ _03899_ _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10128__I _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11401__A2 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10332_ _04085_ _04087_ _04090_ _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10263_ net109 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10194_ _03940_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05919__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08333__A2 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06344__A1 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10979__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10979__B2 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06647__A2 _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09099__I _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 a_operand[16] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput23 a_operand[26] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput34 a_operand[36] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput45 a_operand[46] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput56 a_operand[56] net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput67 a_operand[8] net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput78 b_operand[18] net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput89 b_operand[28] net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08731__I _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07072__A2 _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09349__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09349__B2 _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07347__I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08021__B2 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10903__A1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ _00808_ _00909_ _00944_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08790_ _02321_ _02329_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07741_ _00818_ _00901_ _01137_ _00902_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07672_ _01199_ _00816_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06335__A1 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09411_ _03085_ _03088_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06623_ _00075_ _00079_ _00153_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09342_ _02339_ _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06350__A4 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06554_ _00017_ _00084_ _00085_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07835__A1 _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09273_ _02665_ _02937_ _02325_ _02938_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__06638__A2 _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06485_ _03444_ _03182_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08224_ _01748_ _01752_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09588__A1 _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08155_ _01628_ _01722_ _01724_ _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11395__A1 _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07106_ _00533_ _00534_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08641__I _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08086_ _01644_ _01646_ _01649_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07063__A2 _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07037_ _00560_ _00563_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06810__A2 _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07257__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06161__I _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09355__A4 _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08988_ _02404_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06574__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10370__A2 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output134_I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07939_ _01416_ _05169_ _01379_ _01484_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_56_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10950_ net30 _03851_ _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09609_ _03202_ _03206_ _03200_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10881_ _04616_ _04683_ _04684_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_44_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09276__B1 _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08816__I _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09579__A1 _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09043__A3 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08251__A1 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11364_ _05206_ _05209_ _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10315_ _04058_ _04064_ _04067_ _04073_ net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__06801__A2 _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11295_ _05052_ _05110_ _05134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10246_ _03989_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08003__A1 _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10177_ _03919_ _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09503__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10321__I _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09806__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07817__A1 _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06270_ _05476_ _05480_ _05481_ _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08490__A1 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08242__A1 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09960_ _03534_ _03686_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08911_ _02545_ _01257_ _02546_ _02547_ _00968_ _02238_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_69_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09891_ _03609_ _03537_ _03611_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08545__A2 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09742__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08842_ _02231_ _02472_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06556__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10352__A2 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08773_ _02395_ _02396_ _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05985_ _01836_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07724_ _05504_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11301__A1 _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07655_ _01153_ _01114_ _01180_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_65_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06606_ _01488_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07586_ _01094_ _01106_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09325_ _02627_ _02693_ _02922_ _02994_ _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06537_ _00001_ _00026_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07808__A1 _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10407__A3 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09256_ _02347_ _02363_ _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input95_I b_operand[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06468_ _05617_ _00000_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08207_ _01703_ _01708_ _01780_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09187_ _02770_ _02787_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06399_ _05608_ _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11368__A1 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08138_ _01538_ _01706_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08233__A1 _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07036__A2 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09981__A1 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08069_ _01554_ _01631_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_134_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10100_ _03829_ _03838_ net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11080_ net107 net32 _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10031_ _02435_ _02336_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10141__I _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10933_ _03832_ _04009_ _04676_ _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10864_ _04591_ _04630_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _04581_ _04590_ _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06066__I _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09016__A3 _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09377__I _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11416_ _05070_ _05264_ _05265_ _05163_ _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08224__A1 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10031__A1 _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11347_ _03861_ _04237_ _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09972__A1 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10582__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06015__B _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11278_ _04937_ _05114_ _05116_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08527__A2 _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10229_ _03930_ _03973_ _03974_ _03979_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_79_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06538__A1 _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05770_ net26 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10098__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07440_ _00855_ _00865_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07371_ net129 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09110_ _02415_ _02642_ _02761_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06322_ _05527_ _05531_ _05292_ _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09041_ _02616_ _02617_ _02369_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06253_ _05421_ _05463_ _05464_ _05465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08215__A1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07018__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06704__I _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06184_ _02737_ _03346_ _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06226__B1 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10226__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09943_ _03577_ _03590_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09715__A1 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09874_ _03409_ _03592_ _03535_ _03533_ _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_58_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10325__A2 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08825_ _02453_ _02414_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_97_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08756_ _02372_ _02377_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05968_ _04247_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input10_I a_operand[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10896__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07707_ _00953_ _00812_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08687_ _02301_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05899_ _03411_ _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07638_ _00877_ _00845_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ _01088_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09246__A3 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ _05104_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10580_ _04357_ _04358_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _02842_ _02848_ _02901_ _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08206__A1 _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11201_ _04842_ _05026_ _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10136__I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06768__A1 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11132_ _04912_ _04956_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08509__A2 _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09706__A1 _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11063_ _04393_ _04235_ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10014_ _03664_ _03743_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05743__A2 _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10916_ _04040_ _04041_ _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07496__A2 _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11029__B1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10847_ _04643_ _04645_ _04646_ _04647_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10778_ _04570_ _04572_ _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10004__A1 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06759__A1 _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06940_ _00466_ _00467_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05982__A2 _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I Operation[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06871_ _03878_ _05280_ _00396_ _05282_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07184__A1 _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08610_ net47 _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05822_ _02661_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09590_ _03177_ _03282_ _03283_ _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06931__A1 _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08541_ _01980_ _02045_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05753_ _01596_ _01662_ _01738_ _01781_ _01141_ _01912_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_54_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08472_ _02067_ _02068_ _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05684_ net1 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07423_ _00943_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10491__A1 _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ net113 _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08436__A1 _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10243__A1 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06305_ _05436_ _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08987__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07285_ _00804_ _00807_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06998__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09024_ _02653_ _02654_ _02668_ _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06236_ _05447_ _02607_ _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06434__I _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09936__A1 _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06167_ _02650_ _02694_ _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10546__A2 _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input58_I a_operand[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06098_ _05296_ _05312_ _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_49_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09926_ _03648_ _03649_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09164__A2 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09857_ _03416_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08808_ _02431_ _02435_ _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08911__A2 _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09788_ _02890_ _02322_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08739_ _02359_ _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11274__A3 _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10701_ _03870_ _03874_ _04488_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10632_ _04316_ _04347_ _04386_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10563_ _04281_ _04324_ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06989__A1 _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10494_ _03910_ _03917_ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11115_ _04873_ _04920_ _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11046_ _04787_ _04790_ _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09155__A2 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07469__A2 _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10473__A1 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08418__A1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07070_ _00594_ _00595_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06021_ _04822_ _02932_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10528__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07972_ _01377_ _01525_ _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05955__A2 _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09711_ _02513_ _02266_ net62 _02794_ _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_06923_ _00375_ _00380_ _00450_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09642_ _03339_ _03340_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06854_ _00359_ _00382_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_95_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05805_ _02478_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09573_ _03263_ _03264_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06785_ _04691_ _00313_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input112_I b_operand[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08524_ _00770_ _00837_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05736_ _01727_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_64_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10464__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08455_ _02046_ _02050_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06132__A2 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07406_ _00776_ _00928_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08386_ _01904_ _01905_ _01974_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08644__I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07337_ _00847_ _00852_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05891__A1 _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09082__A1 _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07268_ _00790_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09007_ _02603_ _02599_ _02602_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06219_ _05377_ _05382_ _05393_ _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07199_ _00722_ _00723_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10519__A2 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09385__A2 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output164_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05946__A2 _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09137__A2 _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09909_ _03605_ _03631_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07723__I _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10615_ _03880_ _04335_ _01123_ _04396_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10546_ _04316_ _04317_ _04321_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07623__A2 _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10477_ _04242_ _04243_ _04246_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11029_ _03857_ _01858_ _04065_ _04626_ _04817_ _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__08729__I _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10694__A1 _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06570_ _02313_ _01531_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09300__A2 _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _01809_ _01817_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06185__S _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06665__A3 _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08171_ _00789_ _01223_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10749__A2 _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07122_ _00541_ _00547_ _00647_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__A1 _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07053_ _00319_ _00579_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06004_ _02791_ _04637_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput133 net133 ALU_Output[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput144 net144 ALU_Output[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput155 net155 ALU_Output[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07378__A1 _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput166 net166 ALU_Output[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput177 net177 ALU_Output[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput188 net188 ALU_Output[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput199 net199 Exception[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10382__B1 _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07955_ _01502_ _01506_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06906_ _00336_ _00385_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08639__I _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07886_ _01365_ _01399_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09625_ _03319_ _03320_ _03321_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10685__A1 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06837_ _03640_ _05365_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10685__B2 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07550__A1 _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07550__B2 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09556_ _03227_ _03245_ _03246_ _01976_ _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06768_ _03564_ _02704_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08507_ _02002_ _02005_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05719_ _01542_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09487_ _03103_ _03107_ _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06699_ _00218_ _00208_ _00222_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10988__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08438_ _00918_ _00890_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09055__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11014__B _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08369_ _01951_ _01957_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10400_ _04149_ _04151_ _04164_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_11380_ _05173_ _05177_ _05226_ _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10853__B _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10331_ _04085_ _04087_ _04090_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10262_ _03858_ _04014_ _04015_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09358__A2 _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10144__I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10193_ _03939_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06041__A1 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06344__A2 _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10979__A2 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput13 a_operand[17] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput24 a_operand[27] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput35 a_operand[37] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput46 a_operand[47] net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput57 a_operand[57] net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput68 a_operand[9] net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10600__A1 _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput79 b_operand[19] net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10529_ _03818_ _04237_ _04195_ _03811_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09349__A2 _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08021__A2 _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07740_ _00902_ _01203_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07363__I _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10667__A1 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07671_ _01188_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07532__A1 _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09410_ _02923_ _03086_ _03016_ _03087_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_53_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06622_ _01770_ _02291_ _00080_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ _03009_ _03012_ _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06553_ _00020_ _00022_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06099__A1 _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09272_ _02476_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06707__I _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06484_ _00014_ _00015_ _00016_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_33_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08223_ _01796_ _01797_ _01798_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08154_ _01561_ _01723_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07599__A1 _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11395__A2 _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07105_ _00491_ _00630_ _00544_ _00545_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08085_ _01191_ _01647_ _01648_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06271__A1 _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07036_ _02269_ _02704_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input40_I a_operand[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08987_ _01118_ _02620_ _02623_ _02628_ _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07771__A1 _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06574__A2 _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07771__B2 _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07938_ _01489_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07273__I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10658__A1 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07869_ _01256_ _01410_ _01414_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09608_ _03200_ _03202_ _03206_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_43_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10880_ _04191_ _04005_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09539_ _03227_ _03142_ _03228_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08079__A2 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09276__A1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09276__B2 _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07826__A2 _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10139__I _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09579__A2 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08832__I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11386__A2 _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11363_ _05041_ _05207_ _05208_ _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08251__A2 _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06262__A1 _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10314_ _04060_ _00421_ _04068_ _04604_ _04072_ _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_11294_ _05054_ _05109_ _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11138__A2 _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10245_ _03996_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08003__A2 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09200__A1 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10176_ _03919_ _03920_ _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10897__A1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06565__A2 _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07762__A1 _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10649__A1 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11074__A1 _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05828__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10821__A1 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09019__A1 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08742__I _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07358__I _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08910_ _02524_ _02545_ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09890_ _03532_ _03610_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06005__A1 _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09742__A2 _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08841_ _02471_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06556__A2 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08772_ _02394_ _02376_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05984_ _04410_ _04420_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07723_ _00905_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07654_ _01153_ _01114_ _01180_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_53_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06605_ _05446_ _00060_ _00122_ _05496_ _00136_ net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__09258__A1 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07585_ _01101_ _01105_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11065__A1 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09324_ _02920_ _02923_ _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11065__B2 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06536_ _00028_ _00066_ _00067_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09255_ _02916_ _02917_ _02918_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06467_ _05619_ _05632_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08481__A2 _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08206_ _00757_ _00775_ _01709_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input88_I b_operand[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08652__I _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06398_ _05547_ _05606_ _05607_ _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09186_ net117 _02373_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08137_ _00918_ _00833_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08233__A2 _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07268__I _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08068_ _01625_ _01628_ _01630_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09981__A2 _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07019_ _00544_ _00545_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10030_ _02278_ _02327_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10879__A1 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09733__A2 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07744__A1 _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09497__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10932_ _04664_ _04718_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10863_ _04592_ _04629_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10794_ _04585_ _04589_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06483__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09016__A4 _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11415_ _05162_ _05164_ _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10031__A2 _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11346_ _05187_ _05189_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07983__A1 _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06786__A2 _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11277_ _05113_ _05012_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10228_ _03975_ _03978_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07735__A1 _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10159_ _03902_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10098__A2 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08160__A1 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06171__B1 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07370_ _00892_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06321_ _05527_ _05531_ _05532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06252_ _05420_ _05423_ _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09040_ _01430_ _02686_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06474__A1 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10270__A2 _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06183_ _03313_ _05339_ _05395_ _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09412__A1 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10558__B1 _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06226__A1 _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06226__B2 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09942_ _03665_ _03666_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09715__A2 _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09873_ _03114_ _02656_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07726__A1 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10242__I _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ _02336_ _02452_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08755_ _02376_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09479__A1 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05967_ _04236_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07706_ _01214_ _01220_ _01236_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_72_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08686_ _02300_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07551__I _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05898_ _03487_ _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07637_ _01096_ _01161_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07568_ net27 _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09307_ _02812_ _02956_ _02969_ _02975_ net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06519_ _03629_ _03661_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07499_ _00998_ _01019_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06465__A1 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09238_ _02778_ _02789_ _02847_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07662__B1 _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10261__A2 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output194_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11022__B _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10417__I _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08206__A2 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09169_ _00137_ _02763_ _02811_ _02812_ _02826_ net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_107_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11200_ _04756_ _05031_ _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06768__A2 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11131_ _04332_ _04908_ _04913_ _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_107_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11062_ _04879_ _04881_ _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_49_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07717__A1 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10013_ _03664_ _03743_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10152__I _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__A1 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ _04049_ _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09890__A1 _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11029__A1 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11029__B2 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06077__I _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _04552_ _02822_ _05585_ _04559_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10777_ _04500_ _04543_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10327__I _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10004__A2 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11329_ _05068_ _05072_ _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10960__B1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _02063_ _00130_ _00394_ _00210_ _00398_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_95_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07184__A2 _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05821_ _02650_ _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08540_ _01980_ _02045_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05752_ _01825_ _01901_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07371__I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A1 _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08471_ _01986_ _02044_ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05683_ net3 _01151_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09881__A1 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07422_ _00944_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07353_ _00873_ _00875_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08436__A2 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06304_ _05509_ _05511_ _05512_ _05515_ _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06447__B2 _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07284_ _00806_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09023_ _02662_ _02664_ _02667_ _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10237__I _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06235_ _02564_ _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09936__A2 _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06166_ _01868_ _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06097_ _05297_ _05299_ _05311_ _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_49_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09925_ _03552_ _03558_ _03551_ _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_59_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09856_ _03526_ _03538_ _03572_ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07175__A2 _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08807_ _02433_ _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09787_ _02818_ _03393_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06999_ _00363_ _00477_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11259__A1 _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08738_ _02358_ _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08669_ _02282_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output207_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _03876_ _03885_ _04480_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10631_ _04316_ _04347_ _04386_ _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_41_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08427__A2 _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09624__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10562_ _00137_ _04277_ _04325_ _02812_ _04339_ net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_10_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10147__I _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10493_ _04027_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07650__A3 _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11114_ _04861_ _04866_ _04936_ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11045_ _04703_ _04862_ _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05704__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09863__B2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10473__A2 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07874__B1 _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10829_ _04594_ _04611_ _04628_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_60_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06020_ _01270_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09379__B1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09918__A2 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08750__I _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07366__I _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06062__C1 _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ _00903_ _01085_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09710_ _03414_ _03328_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06922_ _00377_ _00449_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08354__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09641_ _03259_ _03214_ _03338_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06853_ _00371_ _00381_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05804_ net85 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09572_ _03168_ _03211_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06784_ _03835_ _00224_ _02161_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08106__A1 _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08106__B2 _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08523_ net10 _00837_ _00852_ _00770_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05735_ _01683_ _01716_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input105_I b_operand[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10464__A2 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08454_ _01893_ _02048_ _02049_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07405_ _00778_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08385_ _01899_ _01903_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_50_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07336_ _00858_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05891__A2 _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07267_ _00789_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input70_I b_operand[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09006_ _02593_ _02648_ _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08660__I _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06218_ _01412_ _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07198_ _00652_ _00659_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06149_ _05300_ _02715_ _03269_ _01553_ _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_132_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07276__I _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08593__A1 _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output157_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09908_ _03608_ _03630_ _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09839_ _03436_ _03437_ _03435_ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__B1 _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09845__A1 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10586__B _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11404__A1 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10614_ _00418_ _04395_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10545_ _04318_ _04320_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_41_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06831__A1 _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10476_ _04081_ _04127_ _04244_ _04245_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__08584__A1 _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10391__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__A1 _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11028_ _04834_ _04844_ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06898__A1 _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07862__A3 _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08170_ _00780_ _00765_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06265__I _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07121_ _00543_ _00546_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07075__A1 _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08811__A2 _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07052_ _00427_ _00502_ _00578_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06003_ _01640_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput134 net134 ALU_Output[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput145 net145 ALU_Output[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput156 net156 ALU_Output[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07378__A2 _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput167 net167 ALU_Output[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput178 net178 ALU_Output[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10382__A1 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput189 net189 ALU_Output[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10382__B2 _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07954_ _00925_ _00946_ _01505_ _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08327__A1 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06905_ _00340_ _00384_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07885_ _01365_ _01399_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09624_ _02671_ _02272_ _03236_ _02234_ _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06836_ _00361_ _00362_ _00364_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10685__A2 _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07550__A2 _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09555_ _03227_ _03245_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06767_ _02368_ _03258_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08506_ _02003_ _02004_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05718_ _01531_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09486_ _03110_ _03130_ _03169_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06698_ _00218_ _00208_ _00222_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08437_ _02028_ _02030_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08368_ _00906_ _00809_ _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07319_ _00830_ _00835_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08299_ _00418_ _00771_ _00940_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10330_ _04074_ _04089_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10425__I _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10261_ _03853_ _03857_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08566__A1 _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10192_ _03938_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06041__A2 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10160__I _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09818__A1 _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06085__I _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 a_operand[18] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput25 a_operand[28] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput36 a_operand[38] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput47 a_operand[48] net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput58 a_operand[58] net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10528_ _03897_ _03809_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10600__A2 _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput69 b_operand[0] net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10459_ _03913_ _03841_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10667__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07670_ _01149_ _01150_ _01198_ net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07532__A2 _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06621_ _00068_ _00150_ _00151_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09340_ _03005_ _03010_ _03011_ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10419__A2 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06552_ _00020_ _00022_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09271_ _02312_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11092__A2 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06483_ net21 _02943_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08222_ _01713_ _01734_ _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08153_ _00797_ net49 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08796__A1 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07104_ _02423_ _03564_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08084_ _00810_ _01381_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07035_ _02172_ _05324_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06271__A2 _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10355__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06559__B1 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08986_ _02624_ _05280_ _05507_ _02542_ _02627_ _01577_ _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_102_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input33_I a_operand[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07554__I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07771__A2 _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07937_ _00791_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07868_ _01879_ _01413_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__A2 _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09607_ _03285_ _03301_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06819_ _00330_ _00347_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07799_ _01256_ _05169_ _01379_ _01273_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ _02458_ _02459_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09276__A2 _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09469_ _04930_ _03072_ _03140_ _03152_ net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09028__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11362_ _05045_ _05111_ _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10313_ _00951_ _04069_ _04071_ _00959_ _04070_ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__10155__I _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06262__A2 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11293_ _05048_ _05051_ _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10244_ _03993_ _03995_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10346__A1 _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07211__A1 _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10175_ net34 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10897__A2 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07762__A2 _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06565__A3 _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10649__A2 _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07278__A1 _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11074__A2 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05828__A2 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10821__A2 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09019__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08778__A1 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10585__A1 _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10337__A1 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ _02447_ _02470_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06005__A2 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10888__A2 _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07753__A2 _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _02394_ _02376_ _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05983_ _04118_ _04182_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07722_ _05502_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07653_ _01154_ _01179_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_81_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06604_ _02335_ _05644_ _00125_ _05648_ _00135_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_25_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07584_ _01090_ _01103_ _01104_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09258__A2 _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09323_ _02919_ _02933_ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06535_ _00027_ _00031_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _02784_ _02861_ _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06466_ _05673_ _05638_ _05674_ _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08205_ _01698_ _01758_ _01778_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09185_ _02778_ _02789_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06397_ _05543_ _05485_ _05550_ _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08136_ _01612_ _01642_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10576__A1 _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08067_ _00906_ _01074_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07018_ _02368_ _02586_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10879__A2 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07284__I _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08969_ _02520_ _02576_ _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10931_ _04667_ _04717_ _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10862_ _04585_ _04589_ _04663_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06180__A1 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _04523_ _04586_ _04588_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10803__A2 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06483__A2 _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11414_ _04005_ _03904_ _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11345_ _05095_ _05188_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07983__A2 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10319__A1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11276_ _05113_ _05012_ _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10613__I _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10227_ _03976_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10158_ net36 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10089_ _03826_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06171__A1 _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06171__B2 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06320_ _02629_ _05528_ _05529_ _05530_ _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08753__I _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06251_ _05420_ _05423_ _05463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06474__A2 _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07369__I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06182_ _05318_ _03302_ _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10558__B2 _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06226__A2 _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09941_ _03605_ _03631_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09176__A1 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10523__I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09872_ _03577_ _03590_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07726__A2 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08923__A1 _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _02340_ _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08754_ _02375_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05966_ _01336_ _04065_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09479__A2 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07705_ _01235_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08685_ _02299_ _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05897_ _03378_ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07636_ _00749_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06162__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07567_ _01085_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11038__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06892__B _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09100__A1 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09306_ _02957_ _02973_ _02974_ _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06518_ _00048_ _05435_ _03672_ _05437_ _00050_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07498_ _01016_ _01018_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_139_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10797__A1 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09237_ _02839_ _02879_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07662__A1 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06449_ _02445_ _03618_ _05658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09168_ _02321_ _02744_ _02816_ _02751_ _02825_ _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__10549__A1 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output187_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08119_ _01685_ _01651_ _00126_ _01579_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11210__A2 _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09099_ _04075_ _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11130_ _04882_ _04890_ _04954_ _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07965__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05976__A1 _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11061_ _04862_ _04880_ _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10012_ _03731_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08914__A1 _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10914_ _04659_ _04720_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06153__A1 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10845_ _04040_ _04552_ _01193_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11029__A2 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10776_ _04503_ _04542_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10788__A1 _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06208__A2 _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11328_ _05069_ _05070_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10960__A1 _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10960__B2 _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11259_ _04960_ _05095_ _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07708__A2 _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08905__A1 _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10712__A1 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05820_ _02639_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08748__I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10499__B _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05751_ _01781_ _01890_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08133__A2 _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ _01989_ _02043_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06144__A1 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05682_ net4 _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10011__C _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07421_ _00943_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__A1 _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07352_ _00874_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09633__A2 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06303_ _05514_ _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06447__A2 _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07283_ _00805_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09022_ _02665_ _02655_ _02560_ _02666_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_06234_ _05445_ _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06165_ _05377_ _05378_ _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06096_ _05306_ _05310_ _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10951__A1 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10253__I _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09924_ _03645_ _03647_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09855_ _03514_ _03525_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_86_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08806_ _02432_ _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09786_ _03493_ _03496_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06998_ _02074_ _01520_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08737_ _02356_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05949_ _01976_ _04043_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06135__A1 _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08668_ _02281_ _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09872__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07619_ _00891_ _00896_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08599_ _02206_ _02207_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10630_ _04342_ _04411_ _04412_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09624__A2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05810__I _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07635__A1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10561_ _03891_ _02744_ _04328_ _02751_ _04338_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_10_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10492_ _03899_ _05498_ _04256_ _05503_ _04263_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_108_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09388__A1 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05949__A1 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _03831_ _04019_ _04867_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10163__I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11044_ _03861_ _04297_ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08363__A2 _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09560__A1 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07571__B1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__A1 _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07874__B2 _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10828_ _04619_ _04627_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_13_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10759_ _04470_ _04279_ _05321_ _04487_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_9_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09379__A1 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09379__B2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08051__A1 _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10933__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06062__B1 _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10073__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07970_ _01453_ _01456_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06062__C2 _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06921_ _05515_ _00373_ _00378_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_68_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08354__A2 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09640_ _03259_ _03214_ _03338_ _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06852_ _00375_ _00380_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05803_ net21 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09571_ _03262_ _03210_ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06783_ _00138_ _00227_ _00312_ net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08106__A2 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08522_ _02012_ _02018_ _02123_ _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05734_ _01607_ _01151_ _01694_ _01705_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_82_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08453_ _02047_ _01967_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07404_ _00783_ _00786_ _00795_ _00925_ _00926_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_11_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08384_ _01869_ _01871_ _01885_ _01973_ net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09102__I _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ _00846_ _00849_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07617__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07266_ net7 _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08941__I _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09005_ _02377_ _02383_ _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06217_ _05394_ _05377_ _05382_ _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07197_ _00654_ _00658_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11177__A1 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input63_I a_operand[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06148_ _05324_ _01553_ _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10924__A1 _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08593__A2 _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06079_ _01694_ _01955_ _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09907_ _03612_ _03628_ _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09838_ _03551_ _03554_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06356__A1 _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07292__I _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05805__I _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09769_ _03475_ _03478_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__A1 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__B2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09012__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10158__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10613_ _04394_ _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10544_ _04228_ _04319_ _04298_ _04201_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_41_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07084__A2 _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08281__A1 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10475_ _04184_ _04201_ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11168__A1 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07467__I _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09781__A1 _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06595__A1 _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10391__A2 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__A2 _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09533__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11027_ _01792_ _04817_ _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10143__A2 _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09631__B _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09297__B1 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07847__A1 _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07120_ _00645_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09857__I _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07051_ _00429_ _00430_ _00501_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11159__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06002_ _04615_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08024__A1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08024__B2 _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput135 net135 ALU_Output[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput146 net146 ALU_Output[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput157 net157 ALU_Output[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09772__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput168 net168 ALU_Output[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput179 net179 ALU_Output[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10382__A2 _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07953_ _01503_ _00943_ _01504_ _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10531__I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06904_ _00329_ _00333_ _00431_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07884_ _05665_ _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11331__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10134__A2 _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09623_ _03236_ _02487_ _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06835_ _00265_ _00363_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09554_ _02428_ _02556_ _03244_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06766_ _00193_ _00294_ _00295_ _00095_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_24_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08505_ _01957_ _02104_ _02015_ _02016_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_52_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05717_ _01520_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09485_ _03112_ _03129_ _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06697_ _00222_ _00226_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08436_ _01916_ _02029_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10842__B1 _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08367_ _00904_ _00813_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07318_ _00831_ _00836_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08671__I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08263__A1 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08298_ _01859_ _01872_ _01193_ _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10070__A1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07249_ net75 _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07287__I _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10260_ _04003_ _04011_ _04013_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08015__A1 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11030__C _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08566__A2 _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10191_ _03937_ _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06577__A1 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11322__A1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08846__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09818__A2 _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 a_operand[19] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput26 a_operand[29] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput37 a_operand[39] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput48 a_operand[49] net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput59 a_operand[59] net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_10527_ _04296_ _04300_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10600__A3 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08006__A1 _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10458_ _04199_ _04202_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10389_ _04115_ _04119_ _04152_ _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06568__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11313__A1 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06050__B _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06620_ _00072_ _00116_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06740__A1 _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07660__I _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09809__A2 _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06551_ _00002_ _00009_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09270_ _02219_ net121 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06482_ net22 net77 _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11092__A3 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08221_ _01754_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08152_ _01625_ _01630_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08245__A1 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09442__B1 _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07103_ _00628_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08083_ _00904_ _00874_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07034_ _00354_ _00560_ _00464_ _00462_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08985_ _02626_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07936_ _00979_ _01486_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11304__A1 _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10107__A2 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input26_I a_operand[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07867_ _01411_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09606_ _03286_ _03300_ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08666__I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06818_ net25 _02943_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07798_ _04323_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06731__A1 _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09537_ _02436_ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06749_ _02478_ _02650_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09468_ _02458_ _01251_ _03144_ _03151_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08419_ _02011_ _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09399_ _02991_ _03075_ _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08236__A1 _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__A1 _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09984__A1 _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11361_ _05045_ _05111_ _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_125_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10312_ _04059_ _04070_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11292_ _05129_ _05130_ _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09736__A1 _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10243_ _03990_ _03994_ _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10174_ net98 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10171__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09503__A4 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07278__A2 _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08227__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10034__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08778__A2 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10585__A2 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10337__A2 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10081__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08770_ _02393_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05982_ _01781_ _01585_ _03128_ _01141_ _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07721_ _01252_ _01253_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07652_ _01176_ _01178_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06713__A1 _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06174__C1 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07390__I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06713__B2 _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05903__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06603_ _00127_ _00128_ _00132_ _00134_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_80_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07583_ _00830_ _00849_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06534_ _00027_ _00031_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09322_ _02316_ _02503_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08466__A1 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06465_ _05556_ _05572_ _05633_ _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09253_ _02784_ _02861_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08204_ _01700_ _01757_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08218__A1 _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09184_ _02342_ _02384_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06396_ _05543_ _05485_ _05550_ _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08135_ _01638_ _01652_ _01702_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10256__I _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08066_ net130 net60 _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09718__A1 _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07017_ _05524_ _00539_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08968_ _02547_ _02608_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07919_ _01373_ _01388_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08899_ _02223_ _02239_ _02254_ _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09497__A3 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10930_ _04659_ _04720_ _04737_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05813__I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10500__A2 _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10861_ _03831_ _04041_ _04590_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06180__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10792_ _04436_ _04587_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09654__B1 _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10016__A1 _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11413_ _05260_ _05261_ _05262_ _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10166__I _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11344_ net46 _03934_ _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07432__A2 _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09709__A1 _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11275_ _04941_ _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10226_ _03928_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10157_ _03899_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06943__A1 _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10088_ net94 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07424__B _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05723__I _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08160__A3 _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06171__A2 _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06250_ _05459_ _05424_ _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10007__A1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10076__I _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06181_ _05393_ _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10558__A2 _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09940_ _03573_ _03604_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09871_ _03583_ _03589_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08822_ _02450_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06934__A1 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08753_ _02374_ _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05965_ _03128_ _04171_ _04182_ _04215_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07704_ _01226_ _01234_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input128_I b_operand[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08684_ _02298_ _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05896_ _03422_ _03465_ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10494__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07635_ _01031_ _01158_ _01159_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07566_ net102 _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09100__A2 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09305_ _02957_ _02973_ _01139_ _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06517_ _05650_ _00049_ _01368_ _00043_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_70_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07497_ _00993_ _01017_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input93_I b_operand[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09236_ _02841_ _02877_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07662__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06448_ _05446_ _05601_ _05643_ _05496_ _05657_ net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__06870__B1 _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09167_ _02821_ _02823_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06379_ _05331_ _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08118_ _00932_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06217__A3 _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09098_ _02747_ _02749_ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08049_ _01535_ _01548_ _01609_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05976__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11060_ net43 _03948_ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07178__A1 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10011_ _03649_ _03740_ _03741_ _03733_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_1_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06925__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10721__A2 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10913_ _04662_ _04719_ _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06153__A2 _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08854__I _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10844_ _04644_ _04334_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11029__A3 _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _04567_ _04568_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__A1 _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11327_ _05002_ _05168_ _05081_ _05083_ _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_141_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05718__I _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10960__A2 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09158__A2 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11258_ net45 _03950_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07169__A1 _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10209_ _03957_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11189_ _04935_ _05018_ _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05750_ _01847_ _01879_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10476__A1 _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05681_ _01130_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07341__A1 _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07420_ _00942_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08764__I _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10228__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07351_ net113 _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10779__A2 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06302_ _05513_ _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07282_ net131 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06284__I _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09021_ _02350_ _02484_ _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06233_ _05444_ _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06164_ _05329_ _05376_ _05337_ _05378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_132_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06095_ _05308_ _05309_ _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10951__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09923_ _03471_ _03545_ _03646_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09854_ _03569_ _03570_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09544__B _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ net61 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09785_ _03494_ _03495_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06997_ _00479_ _00483_ _00523_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08736_ _02355_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05948_ _02042_ _04032_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08667_ _02279_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06135__A2 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05879_ _03248_ _03280_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08674__I _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07618_ _01112_ _01115_ _01133_ _01142_ net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08598_ _02128_ _02136_ _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07549_ _00881_ _00049_ _01368_ _01040_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_139_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10560_ _04333_ _04336_ _04337_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_139_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09219_ _02838_ _02880_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10491_ _01379_ _04253_ _04261_ _04262_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07399__A1 _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08060__A2 _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11112_ _04934_ _04927_ _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11043_ _04783_ _04859_ _04860_ _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08899__A1 _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09560__A2 _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08115__A3 _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__A2 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10827_ _04622_ _04625_ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07626__A2 _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10758_ _04041_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10689_ _03869_ _05498_ _04469_ _05503_ _04476_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09379__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07149__B _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06062__A1 _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10933__A2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06920_ _00349_ _00356_ _00447_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10697__A1 _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06851_ _00377_ _00379_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05802_ _02390_ _02423_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09570_ _03170_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06782_ _00230_ _00236_ _00243_ _00311_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_83_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08521_ _02014_ _02017_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05733_ _01390_ _01184_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08452_ _02047_ _01967_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05911__I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07403_ _00791_ _00794_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08383_ _00425_ _01972_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07334_ _00742_ _00744_ _00769_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11413__A3 _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07265_ _00783_ _00787_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09004_ _02573_ _02609_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06216_ _05403_ _05428_ _05429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07196_ _00714_ _00717_ _00720_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_117_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10264__I _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06147_ _05359_ _05360_ _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10924__A2 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input56_I a_operand[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ _05287_ _05289_ _05292_ _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09906_ _03617_ _03627_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__I _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09837_ _03552_ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09768_ _03388_ _03477_ _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ net54 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09699_ _03328_ _03329_ _03318_ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06108__A2 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05821__I _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10612_ net103 _04393_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_41_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10612__A1 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10543_ _03927_ _03953_ _03965_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08281__A2 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10474_ _04200_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11168__A2 _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10174__I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06595__A2 _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07483__I _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _03847_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10679__A1 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09297__B2 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09049__A1 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07050_ _00572_ _00576_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11159__A2 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06001_ _01205_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09757__C1 _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08024__A2 _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09221__A1 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10367__B1 _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput136 net136 ALU_Output[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput147 net147 ALU_Output[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput158 net158 ALU_Output[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09772__A2 _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput169 net169 ALU_Output[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08980__B1 _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07952_ _00920_ _00916_ _00802_ _01349_ _00801_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_68_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07393__I _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05906__I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06903_ _01760_ _03856_ _00334_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07883_ _00923_ _01427_ _01428_ _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07535__A1 _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11331__A2 _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ _02221_ _02273_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06834_ net92 net13 _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09553_ _02829_ _02555_ _03243_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06765_ _02543_ _03455_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input110_I b_operand[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08504_ _00799_ _00905_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05716_ net13 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09484_ _03163_ _03167_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06696_ _04951_ _00224_ _00225_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08435_ net10 _00850_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10842__A1 _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10842__B2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ _01719_ _01945_ _01831_ _01828_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07317_ _00839_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09460__A1 _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ _00939_ _01257_ _00584_ _01685_ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06274__A1 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07568__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10070__A2 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07248_ _00770_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _02151_ _02661_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06026__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ net33 _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output162_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07774__A1 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06577__A2 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10722__I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05816__I _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09515__A2 _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07526__A1 _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11086__A1 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07829__A2 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10169__I _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08862__I _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 a_operand[1] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10597__B1 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput27 a_operand[2] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xinput38 a_operand[3] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput49 a_operand[4] net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10526_ _04298_ _04299_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10457_ _04176_ _04207_ _04224_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08006__A2 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09203__A1 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10388_ _04116_ _04117_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07765__A1 _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07517__A1 _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11313__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07517__B2 _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11009_ _03853_ _05498_ _04815_ _05503_ _04824_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_77_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07941__I _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11077__A1 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06550_ _00010_ _00025_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10824__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06481_ net20 net79 _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08220_ _01713_ _01734_ _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08151_ _01714_ _01720_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09442__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07388__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07102_ _00611_ _00627_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08082_ _00896_ _01128_ _01544_ _01645_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_07033_ _03694_ _03400_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07756__A1 _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__A2 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ _02355_ _02625_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10760__B1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07935_ _01408_ _01413_ _01484_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11304__A2 _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07866_ _01335_ _00800_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09605_ _03292_ _03296_ _03299_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_84_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input19_I a_operand[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06817_ net26 _01998_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07797_ _01335_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09536_ _03218_ _03224_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06748_ net84 net19 _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_19_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09467_ _03145_ _03146_ _03148_ _03149_ _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08484__A2 _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06679_ _02118_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06495__A1 _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08418_ _01841_ _02010_ _01958_ _01956_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08682__I _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09398_ _02998_ _03040_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08349_ _01827_ _01832_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08236__A2 _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09433__A1 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07298__I _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11360_ _05132_ _05135_ _05205_ _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09984__A2 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07995__A1 _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10311_ _03961_ _03816_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11291_ _04848_ _05122_ _05123_ _05121_ _05118_ _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_106_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10242_ _03992_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08944__B1 _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10173_ _03910_ _03917_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_120_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08857__I _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11059__A1 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06377__I _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10806__A1 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08632__C1 _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07986__A1 _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10509_ _04223_ _04251_ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08033__S _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07738__A1 _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07202__A3 _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06410__A1 _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05981_ _01792_ _01596_ _02042_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07720_ _01191_ _01186_ _01201_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07671__I _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08163__A1 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07651_ _01093_ _01107_ _01177_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06174__B1 _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06713__A2 _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06174__C2 _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06602_ _00048_ _05319_ _00133_ _00056_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07582_ _01102_ _00764_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09321_ _02913_ _02949_ _02990_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06533_ _00063_ _00064_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__A1 _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06477__A1 _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09252_ _02855_ _02908_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06464_ _05556_ _05572_ _05633_ _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08203_ _01774_ _01776_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08218__A2 _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09183_ _02774_ _02805_ _02840_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06395_ _05602_ _05604_ _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08134_ _01639_ _01650_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07977__A1 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08065_ _01446_ _01625_ _01626_ _01560_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07016_ _00368_ _00533_ _00542_ _00481_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09718__A2 _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08967_ _02589_ _02594_ _02606_ _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06952__A2 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07918_ _00744_ _00919_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11289__A1 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08677__I _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08898_ _02530_ _02533_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07581__I _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07849_ _00953_ _01335_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07901__A1 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10860_ _04576_ _04660_ _04661_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09103__B1 _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09519_ _03202_ _03206_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10791_ net39 net97 _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09654__A1 _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09406__A1 _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11412_ _05064_ _05250_ _05159_ _05156_ _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10016__A2 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07968__A1 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11343_ _04019_ _03934_ _03952_ net46 _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09709__A2 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06640__A1 _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11274_ _05041_ _05045_ _05111_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_140_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10182__I _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10225_ _03925_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10156_ _03898_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10087_ _03821_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08145__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08448__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10989_ _04757_ _04802_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06180_ _03422_ _03465_ _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08081__B1 _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10092__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09870_ _03587_ _03588_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ _02321_ _02328_ _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06934__A2 _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ _02373_ _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05964_ _04204_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07703_ _01230_ _01233_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08683_ net57 _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05895_ _03433_ _03455_ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07634_ _00871_ _00848_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10494__A2 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07565_ _00836_ _00753_ _00859_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08439__A2 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09304_ _02970_ _02972_ _02699_ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06516_ _01216_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07647__B1 _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07496_ _00743_ _00831_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07111__A2 _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _02895_ _02896_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06447_ _02434_ _05644_ _05647_ _05648_ _05656_ _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input86_I b_operand[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09166_ _02754_ _02822_ _05585_ _02451_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06870__A1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06378_ _05510_ _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06870__B2 _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08117_ _00776_ _00234_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10549__A3 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09097_ _02689_ _02746_ _02745_ _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06622__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08048_ _01536_ _01547_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07178__A2 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10010_ _03657_ _03734_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09999_ _03728_ _03729_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06925__A2 _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08127__A1 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05824__I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06689__A1 _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10912_ _04664_ _04718_ _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_17_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10843_ _04048_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10774_ _04545_ _04546_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10177__I _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08850__A2 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08870__I _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11326_ _03868_ _03883_ _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11257_ net46 _03842_ _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10208_ _03956_ _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10173__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11188_ _04935_ _05018_ _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06916__A2 _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10139_ _03880_ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_39_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09866__A1 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10476__A2 _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05680_ _01119_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07877__B1 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07341__A2 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07350_ _00872_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11425__A1 _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06301_ net20 net84 _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10087__I _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07281_ _00803_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09020_ _02513_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06232_ _01477_ _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ _05329_ _05376_ _05336_ _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07396__I _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06604__B2 _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06094_ _01270_ _03215_ _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09922_ _03473_ _03544_ _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09853_ _03510_ _03540_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10703__A3 _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ _02430_ _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09784_ _03287_ _03387_ _02358_ _02279_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06996_ _00364_ _00478_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07580__A2 _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08735_ net116 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08020__I _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05947_ _01314_ _04010_ _04021_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ net59 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05878_ _03204_ _03269_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07617_ _01120_ _01138_ _01140_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08597_ _02131_ _02135_ _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11416__A1 _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07548_ _00822_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07096__A1 _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07479_ _00958_ _00999_ _01000_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_139_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09218_ _02839_ _02879_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__I _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output192_I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10490_ _04218_ _02822_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09149_ _02777_ _02804_ _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_135_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07399__A2 _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05819__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11111_ _04853_ _04924_ _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09735__B _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09545__B1 _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11042_ _04786_ _04799_ _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07556__C1 _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08899__A2 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09026__I _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10826_ _04620_ _04623_ _04624_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__11407__A1 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10757_ _04548_ _04549_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10091__B1 _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06834__A1 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10091__C2 _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10688_ _04474_ _04475_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08587__A1 _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05729__I _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09784__B1 _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10394__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11309_ _05148_ _05149_ _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06062__A2 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09645__B _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08339__A1 _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11343__B1 _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06850_ _05513_ _00373_ _00378_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_95_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05801_ _02390_ _02434_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06781_ _00244_ _00310_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08520_ _02121_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05732_ _01455_ net2 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08511__A1 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08451_ _01896_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07402_ _00801_ _00910_ _00923_ _00924_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_23_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08382_ _01888_ _01971_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07333_ _00855_ _00768_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08814__A2 _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06825__A1 _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07264_ _00786_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09003_ _02610_ _02609_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06215_ _05405_ _05427_ _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07195_ _00710_ _00718_ _00719_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08578__A1 _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06146_ net82 _05360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10385__A1 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07250__A1 _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06077_ _05291_ _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input49_I a_operand[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09905_ _03626_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11376__I _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07002__A1 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09836_ _03547_ _03550_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09767_ _03386_ _03391_ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06979_ _00404_ _00406_ _00424_ _00506_ net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08718_ _02336_ _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _03384_ _03401_ _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_27_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output205_I net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08649_ _02259_ _02260_ _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10611_ net39 _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10542_ _04227_ _04240_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10473_ _03943_ _03905_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10376__A1 _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07792__A2 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10190__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11025_ _04018_ _04171_ _04840_ _04215_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10679__A2 _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__A2 _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10851__A2 _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09049__A2 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10809_ _03902_ _03907_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10365__I _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06000_ _04593_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09757__B1 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09757__C2 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10367__A1 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10367__B2 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput137 net137 ALU_Output[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput148 net148 ALU_Output[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09375__B _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput159 net159 ALU_Output[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08980__A1 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07951_ _01416_ _00916_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08980__B2 _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06902_ _00324_ _00387_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07882_ _00923_ _01427_ _05445_ _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09621_ _03188_ _03201_ _03304_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06833_ _02151_ _05413_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09552_ _02284_ _03069_ _02427_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06764_ _03465_ _00194_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08503_ _02102_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05715_ _01292_ _01314_ _01498_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09483_ _03164_ _03166_ _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06695_ _02258_ _03813_ _04691_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08434_ net11 _00767_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input103_I b_operand[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10842__A2 _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08365_ _01730_ _01951_ _01952_ _01261_ _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_134_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07316_ _00832_ _00838_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08296_ _01008_ _01875_ _01877_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09460__A2 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07247_ net11 _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07178_ _03694_ _02500_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06129_ _05337_ _05341_ _05342_ _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07774__A2 _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07517__C _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09819_ _02285_ _02656_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10530__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09279__A2 _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05832__I _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11086__A2 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10597__A1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 a_operand[20] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput28 a_operand[30] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10597__B2 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10525_ _03913_ _03949_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10185__I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput39 a_operand[40] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09739__B1 _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10456_ _04178_ _04206_ _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06017__A2 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11010__A2 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10387_ _04101_ _04120_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07765__A2 _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11008_ _04820_ _04821_ _04823_ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05742__I _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10824__A2 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06480_ _05555_ _05616_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09690__A2 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08150_ _01715_ _01717_ _01719_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07101_ _00626_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10095__I _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08081_ _00895_ _00820_ _01381_ _00893_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07032_ _00556_ _00558_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07205__A1 _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05917__I _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ net52 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10760__B2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07934_ _01484_ _01408_ _01413_ _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07865_ _05506_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09604_ _03293_ _03297_ _03298_ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06816_ _00275_ _00281_ _00344_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07796_ _01334_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09535_ _03222_ _03223_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06747_ _00100_ _00266_ _00276_ _00170_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09130__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09466_ _03053_ _05437_ _01189_ _03067_ _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10815__A2 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06678_ _00207_ _00208_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06495__A2 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07692__A1 _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ _00798_ _00809_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09397_ _02982_ _03046_ _03044_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08348_ _01827_ _01832_ _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09433__A2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08279_ _01767_ _01860_ _05245_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10310_ _03836_ _04060_ _03817_ _03832_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07995__A2 _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11290_ _05112_ _05117_ _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09197__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10241_ _03990_ _03992_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08944__A1 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10172_ _03916_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08944__B2 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11059__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09121__A1 _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10806__A2 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09672__A2 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06486__A2 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07435__A1 _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11231__A2 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08632__B1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07986__A2 _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10508_ _04280_ _04250_ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10439_ _04178_ _04206_ _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_98_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05737__I _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08935__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05980_ _04377_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09360__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07650_ _00755_ _00821_ _01091_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06174__A1 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06174__B2 _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06601_ _05518_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07910__A2 _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07581_ _01074_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05921__A1 _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09320_ _02915_ _02948_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06532_ _05672_ _00034_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__A2 _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07123__B1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09251_ _02863_ _02874_ _02914_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06463_ _05635_ _05670_ _05671_ _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08202_ _01692_ _01761_ _01775_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09182_ _02777_ _02804_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06394_ _05542_ _05603_ _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08133_ _00954_ _00774_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09966__A3 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08064_ _01557_ _01561_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07015_ _00480_ _00482_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10733__A1 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08966_ _02604_ _02605_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input31_I a_operand[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07917_ _01449_ _01465_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08897_ _05445_ _02531_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08154__A2 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ _01366_ _01391_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07779_ _01313_ _01316_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09103__B2 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09518_ _03121_ _03203_ _03205_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10790_ _04522_ _04524_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09654__A2 _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ _03110_ _03130_ _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11411_ _03860_ _03894_ _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09738__B _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11342_ _05078_ _05085_ _05185_ _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08090__A1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11273_ _05052_ _05110_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06640__A2 _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10224_ _03909_ _03916_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_121_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10155_ _03897_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10086_ _03821_ _03822_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_94_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10488__B1 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09893__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10988_ _04759_ _04779_ _04801_ _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_90_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07947__I _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08081__A1 _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08081__B2 _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08820_ _02369_ _02448_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08751_ net51 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05963_ _04193_ _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07702_ _01228_ _01231_ _01232_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08682_ _02296_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05894_ _03444_ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06147__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07633_ _01157_ _00764_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07895__A1 _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07564_ _01055_ _01059_ _01082_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09636__A2 _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09303_ _02317_ _02971_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06515_ _02291_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07647__A1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07495_ _01013_ _01014_ _01015_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09234_ _02835_ _02881_ _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06446_ _05649_ _05654_ _05655_ _05656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08018__I _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09165_ _05436_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06377_ _02379_ _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06870__A2 _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08116_ _00964_ _01681_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input79_I b_operand[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09096_ _02745_ _02689_ _02746_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__10954__A1 _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08047_ _00954_ _00781_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06622__A2 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06386__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _02259_ _02539_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08949_ _00138_ _02558_ _02588_ net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09324__A1 _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11131__A1 _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10911_ _04667_ _04717_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06689__A2 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10842_ _03863_ _01257_ _00968_ _04470_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07638__A1 _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10773_ _04566_ _04544_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11198__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08063__A1 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08602__A3 _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10193__I _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11325_ _05153_ _05166_ _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11256_ _05090_ _05091_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10207_ net32 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11187_ _05013_ _05016_ _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10173__A2 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11370__A1 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10138_ _03879_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10069_ _03746_ _03751_ _03805_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06129__A1 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09866__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07877__A1 _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07877__B2 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08547__B _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09618__A2 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11425__A2 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06300_ _05281_ _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07280_ net67 _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06301__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06231_ _05399_ _05400_ _05443_ net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08054__A1 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06162_ _03084_ _05314_ _05286_ _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06604__A2 _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06093_ _04789_ _05303_ _05307_ _05006_ _05308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09921_ _03565_ _03644_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08357__A2 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__A1 _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09852_ _03512_ _03539_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07626__B _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06368__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05925__I _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08803_ _02429_ _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09783_ _03119_ _03120_ _02345_ _02356_ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06995_ _00485_ _00495_ _00521_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08734_ _02349_ _02353_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05946_ _01260_ _01781_ _03999_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11113__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07868__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08665_ _02277_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05877_ _03258_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07616_ _01120_ _01138_ _01139_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09609__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08596_ _02197_ _02200_ _02203_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07547_ _01065_ _01066_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07478_ _00996_ _00997_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07096__A2 _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09217_ _02841_ _02877_ _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06429_ _05613_ _05633_ _05638_ _05639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08045__A1 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09148_ _02790_ _02803_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_output185_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10927__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10927__B2 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09079_ _02228_ _02341_ _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11110_ _04839_ _04841_ _04847_ _04933_ net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11041_ _04786_ _04799_ _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09545__A1 _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09545__B2 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06359__A1 _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05835__I _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07556__B1 _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07556__C2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07020__A2 _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09848__A2 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10825_ _03877_ _03938_ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10188__I _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11407__A2 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10756_ _04468_ _04472_ _04047_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10091__A1 _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10091__B2 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06834__A2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10687_ _04400_ _01265_ _05585_ _04466_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09784__A1 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11308_ _05075_ _05086_ _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08339__A2 _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11239_ _05067_ _05073_ _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11343__A1 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11343__B2 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05800_ _02423_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06780_ _00246_ _00309_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05731_ _01325_ _01673_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ _01975_ _01980_ _02045_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_63_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06522__A1 _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07401_ _00912_ _00921_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08381_ _01969_ _01970_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07332_ _00763_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07078__A2 _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ _00785_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06825__A2 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06214_ _05419_ _05424_ _05426_ _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09002_ _02637_ _02643_ _02644_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07194_ _02280_ _02596_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09775__A1 _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08578__A2 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06145_ _01086_ _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07250__A2 _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _01966_ _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09904_ _03621_ _03625_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09835_ _03547_ _03550_ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07002__A2 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09766_ _03384_ _03401_ _03474_ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06978_ _00425_ _00505_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06761__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07870__I _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08717_ _02334_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05929_ _02129_ _03824_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09697_ _03385_ _03399_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08648_ net128 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07710__B1 _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08579_ _00772_ _00831_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10610_ _00964_ _04391_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10541_ _03827_ _03894_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10472_ _04189_ _04203_ _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09766__A1 _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08569__A2 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09518__A1 _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11024_ _04018_ _04816_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10808_ _04329_ _04306_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10739_ _04217_ _04526_ _04530_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_126_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09757__B2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09221__A3 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10367__A2 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput138 net138 ALU_Output[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput149 net149 ALU_Output[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09509__A1 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ _00795_ _01501_ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08980__A2 _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11316__A1 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ _00326_ _00386_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07881_ _01424_ _00945_ _01426_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09620_ _03311_ _03316_ _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06832_ _05359_ _03867_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07940__B1 _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09551_ _03229_ _03231_ _03241_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06763_ _00290_ _00292_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08502_ _02086_ _02101_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05714_ _01379_ _01423_ _01488_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_24_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09482_ _03015_ _03165_ _03099_ _03097_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06694_ _00223_ _00142_ _03803_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08433_ _02025_ _02026_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08364_ _01835_ _01841_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10055__A1 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _00837_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08295_ _01867_ _00938_ _01876_ _01966_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07246_ _00763_ _00768_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09748__A1 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07177_ _00646_ _00700_ _00701_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input61_I a_operand[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06128_ _05337_ _05341_ _05291_ _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07223__A2 _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10291__I _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06059_ _04366_ _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output148_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09818_ _02296_ _03014_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08696__I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06734__A1 _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10530__A2 _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09749_ _02457_ _03456_ _03457_ _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10046__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10466__I _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10597__A2 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput18 a_operand[21] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10524_ _03920_ _04297_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput29 a_operand[31] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_109_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09739__A1 _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09739__B2 _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10455_ _04180_ _04222_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10349__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10386_ _04099_ _04120_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11297__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06973__A1 _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11007_ _04728_ _05517_ _05520_ _04813_ _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08478__A1 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10037__A1 _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07100_ _00619_ _00625_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08080_ _01643_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07453__A2 _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08650__A1 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07031_ _00453_ _00557_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08982_ _02360_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10760__A2 _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07933_ _00917_ _00922_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__A1 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07864_ _01407_ _01408_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06716__A1 _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05933__I _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09603_ _02319_ _02339_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06815_ _00277_ _00280_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07795_ _01333_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09534_ _03045_ _03135_ _03219_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06746_ _05359_ _02226_ _02313_ _01542_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11068__A3 _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09130__A2 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09465_ _03147_ _00983_ _00234_ _02283_ _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06677_ _00124_ _00206_ _00139_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08416_ _01993_ _02007_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07692__A2 _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09396_ _03067_ _03071_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10028__A1 _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08347_ _01910_ _01914_ _01933_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_20_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08278_ _00213_ _00934_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07229_ _00752_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10240_ _03991_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09197__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10171_ _03915_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08944__A2 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07544__B _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10503__A2 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05843__I _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10267__A1 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07683__A2 _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07435__A2 _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08632__A1 _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08632__B2 _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10507_ _04278_ _04248_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09188__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10438_ _04180_ _04188_ _04205_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_97_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _04080_ _01238_ _04130_ _04131_ _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06174__A2 _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06600_ _00129_ _00130_ _00131_ _02302_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07580_ _01098_ _01099_ _01100_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06531_ _05675_ _00033_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07123__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07123__B2 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09250_ _02792_ _02796_ _02801_ _02873_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06462_ _05561_ _05636_ _05634_ _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07674__A2 _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08201_ _01695_ _01696_ _01759_ _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06393_ _05540_ _05574_ _05603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09181_ _02353_ _02539_ _02772_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08132_ _01616_ _01655_ _01699_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10430__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08063_ net132 _01029_ _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05928__I _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07014_ _00540_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09179__A2 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10733__A2 _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08965_ _02603_ _02599_ _02602_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_102_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07916_ _01451_ _01464_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08896_ _02400_ _02472_ _02529_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input24_I a_operand[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ _01371_ _01389_ _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08974__I _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07778_ _01075_ _01311_ _01315_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10249__A1 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09517_ _02227_ _02432_ _03119_ _02658_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09103__A2 _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06729_ _00187_ _00256_ _00258_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ _03112_ _03129_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ _03053_ _04334_ _02421_ _05320_ _03054_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11410_ _04017_ _03928_ _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11341_ _05080_ _05084_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10972__A2 _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11272_ _05054_ _05109_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10223_ _03942_ _03969_ _03972_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_106_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10154_ net100 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10085_ net94 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10488__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08884__I _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10987_ _04783_ _04786_ _04799_ _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07105__B2 _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08081__A2 _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10963__A2 _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06919__A1 _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10715__A2 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08750_ _02371_ _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05962_ _01858_ _01705_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07701_ _01095_ _00844_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08681_ _02295_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05893_ net83 _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11140__A2 _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07632_ _01156_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08794__I _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07563_ _00755_ _00872_ _01057_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09636__A3 _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09302_ _02311_ _02817_ _02330_ _02760_ _02416_ _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06514_ _00045_ _00046_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07647__A2 _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07494_ _00739_ _00836_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10651__A1 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09233_ _02838_ _02880_ _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06445_ _05588_ _05517_ _05520_ _05596_ _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09164_ _02817_ _05589_ _05590_ _02413_ _02820_ _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06376_ _02510_ _05583_ _05584_ _05585_ _05586_ _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08115_ _01667_ _01664_ _01675_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_107_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09095_ _02347_ _02351_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08046_ _01529_ _01567_ _01605_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09021__A1 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09997_ _03724_ _03726_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08948_ _01152_ _02577_ _02579_ _02580_ _02587_ _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_29_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09324__A2 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08879_ _02512_ _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07335__A1 _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11131__A2 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10910_ _04677_ _04716_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10841_ _04640_ _04641_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _04497_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07638__A2 _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08835__A1 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10642__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A2 _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08063__A2 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11324_ _05161_ _05165_ _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11255_ _04999_ _05005_ _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08879__I _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10206_ _03953_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11186_ _05014_ _05015_ _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07574__A1 _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10137_ _03877_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10068_ _03754_ _03804_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09931__C _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08523__B1 _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10881__A1 _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08826__A1 _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06301__A2 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06230_ _05295_ _05429_ _05430_ _05433_ _05442_ _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11189__A2 _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06161_ _04075_ _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06092_ _01119_ _02834_ _02976_ _01575_ _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09920_ _03568_ _03643_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07693__I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09851_ _03566_ _03567_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06368__A2 _05578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08802_ net125 _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11361__A2 _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09782_ _02433_ _02371_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06994_ _00471_ _00484_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08733_ _02352_ _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05945_ _03999_ _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11113__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input126_I b_operand[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08664_ net123 _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07868__A2 _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05876_ net81 _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05941__I _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07615_ _05444_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05879__A1 _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08595_ _02186_ _02201_ _02202_ _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08029__I _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07546_ _00843_ _01064_ _01039_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10624__A1 _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09490__A1 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07477_ _00998_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input91_I b_operand[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09216_ _02849_ _02876_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06428_ _05634_ _05635_ _05637_ _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09147_ _02797_ _02775_ _02801_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06359_ _05567_ _05569_ _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09242__A1 _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09078_ _02508_ _02452_ _02363_ _02666_ _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_output178_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ _01587_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08699__I _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09545__A2 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11040_ _04754_ _04803_ _04857_ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07556__A1 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07556__B2 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10824_ _03887_ _04441_ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08808__A1 _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11407__A3 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10615__A1 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10755_ _04487_ _04468_ _04472_ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09481__A1 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10091__A2 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06682__I _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10686_ _04470_ _05511_ _01073_ _04335_ _04473_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09233__A1 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09784__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11307_ _05058_ _05074_ _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11238_ _05068_ _05072_ _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11343__A2 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11169_ _04908_ _04913_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05730_ _01433_ _01151_ _01455_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05761__I _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06522__A2 _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06078__B _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07400_ _00917_ _00922_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_63_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08380_ _01889_ _01891_ _01968_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_07331_ _00847_ _00853_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07262_ _00784_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09001_ _02637_ _02643_ _04756_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06213_ _05357_ _05370_ _05425_ _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09224__A1 _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08027__A2 _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07193_ _03716_ _03574_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11031__A1 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06144_ _05301_ _05305_ _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09775__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06075_ _05287_ _05289_ _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09903_ _03623_ _03624_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07538__A1 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11334__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09834_ _03548_ _03549_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06210__A1 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09765_ _03385_ _03399_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06977_ _00428_ _00504_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06761__A2 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ _02333_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05928_ _02151_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09696_ _03392_ _03398_ _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_39_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08647_ _02255_ _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10845__A1 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05859_ _03041_ _03052_ _03063_ _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06513__A2 _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08982__I _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08578_ _00793_ _00811_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07529_ _01048_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09463__A1 _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06277__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11270__A1 _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10540_ _04289_ _04294_ _04315_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10471_ _04227_ _04240_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09215__A1 _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07777__A1 _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05846__I _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11325__A2 _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11023_ _04834_ _04837_ _04838_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06201__A1 _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11089__B2 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10807_ _04530_ _04602_ _04603_ _04447_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08257__A2 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06268__A1 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11261__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10064__A2 _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10738_ _03902_ _03919_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07465__B1 _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07301__I _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08009__A2 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10669_ _04370_ _04455_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09757__A2 _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput139 net139 ALU_Output[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09509__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11316__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06991__A2 _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ _00320_ _00426_ _00427_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07880_ _00974_ _01425_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08193__A1 _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06831_ _00265_ _00270_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06743__A2 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07940__B2 _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09550_ _03147_ _00966_ _03235_ _03240_ _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06762_ _00257_ _00291_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08501_ _02100_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10827__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05713_ _01477_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09481_ net55 net117 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08496__A2 _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06693_ _00129_ _03792_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08432_ _01953_ _01960_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ _00797_ _00892_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09445__A1 _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06259__A1 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07314_ _00836_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10055__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08294_ _00939_ _00940_ _00938_ _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07245_ _00767_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07176_ _00648_ _00660_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07759__A1 _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ _05339_ _05340_ _04713_ _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input54_I a_operand[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09138__I _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06058_ _05223_ _02813_ _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_120_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09381__B1 _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09920__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09381__C2 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09817_ _03319_ _03521_ _03530_ _03424_ _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_86_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09748_ _02457_ _03456_ _01139_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__A1 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09679_ _03379_ _03380_ _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09684__A1 _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__B1 _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10523_ net97 _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput19 a_operand[22] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_143_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10454_ _04188_ _04205_ _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09739__A2 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10482__I _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08411__A2 _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10385_ _04485_ _04142_ _04147_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08175__A1 _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11006_ _03857_ _01418_ _01410_ _04644_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10809__A1 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11234__A1 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09978__A2 _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07989__A1 _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08650__A2 _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07030_ net28 _02965_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06661__A1 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08981_ _02621_ _00983_ _02365_ _01265_ _02622_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_114_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07932_ _01480_ _01482_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__A2 _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07863_ _01341_ _01331_ _01347_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10341__B _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09602_ _02323_ _02332_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06814_ _00293_ _00341_ _00342_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07794_ net68 _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09533_ _02835_ _02979_ _03219_ _03221_ _02981_ _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__06110__I _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06745_ _00176_ _00272_ _00274_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08469__A2 _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__A3 _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09464_ _02438_ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06676_ _00140_ _00124_ _00206_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08415_ _02001_ _02006_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09418__A1 _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09395_ _02426_ _02699_ _03070_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08346_ _01920_ _01932_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07429__B1 _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08277_ _00771_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07228_ _00751_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06652__A1 _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07159_ _00639_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10736__B1 _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06404__A1 _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _03914_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output160_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08157__A1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09409__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11216__A1 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10019__A2 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06891__A1 _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__A2 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10506_ _04241_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _04189_ _04203_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_109_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10368_ _03935_ _00240_ _04127_ _01035_ _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07735__B _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10299_ _03846_ _04056_ _04756_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09648__A1 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06530_ _00036_ _00041_ _00061_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08320__A1 _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07123__A2 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08285__C _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06461_ _05561_ _05636_ _05634_ _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_34_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08200_ _01599_ _01659_ _01763_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09180_ _02713_ _02714_ _02836_ _02837_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06392_ _05486_ _05539_ _05574_ _05602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08131_ _01620_ _01654_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06634__A1 _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08062_ _01552_ _01622_ _01623_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_88_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07013_ _00378_ _00539_ _00492_ _00490_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06105__I _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08964_ _02599_ _02602_ _02603_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08139__A1 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07915_ _01452_ _01463_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08895_ _02400_ _02472_ _02529_ _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10071__B _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07846_ _01373_ _01388_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input17_I a_operand[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07777_ _00823_ _01030_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10249__A2 _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09516_ _02793_ net61 net59 _02794_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06728_ _00089_ _00257_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10297__I _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09447_ _03031_ _03118_ _03127_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06659_ _00189_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ _02964_ _04279_ _05321_ _03048_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_138_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08329_ net10 _00766_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11340_ _05182_ _05183_ _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10421__A2 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11271_ _05088_ _05108_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10222_ _03963_ _03965_ _03970_ _03971_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_133_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06928__A2 _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10153_ _03891_ _03895_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10084_ _03820_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09878__A1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10488__A2 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08550__A1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07353__A2 _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10986_ _04791_ _04798_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06864__A1 _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09802__A1 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10176__A1 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07041__A1 _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I a_operand[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05961_ _01585_ _03128_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09869__A1 _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07700_ net113 _01029_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08680_ net121 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05892_ _03356_ _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07631_ net60 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07562_ _01045_ _01046_ _01060_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09097__A2 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09301_ _02317_ _02418_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06513_ _05646_ _05652_ _00043_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07493_ _00846_ _00767_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06304__B1 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09232_ _00762_ _02831_ _02894_ net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06444_ _05650_ _05511_ _05512_ _05653_ _05654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10651__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09163_ _02754_ _04615_ _05591_ _02819_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06375_ _01683_ _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08114_ _01667_ _01664_ _01675_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09094_ _02454_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ _01449_ _01465_ _01566_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07032__A1 _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09996_ _03725_ _03706_ _03616_ _03613_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08947_ _02542_ _01238_ _02583_ _02585_ _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08985__I _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08878_ net111 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11131__A3 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07829_ _01301_ _01370_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_72_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10840_ _04555_ _04549_ _04559_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10771_ _04559_ _04564_ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08835__A2 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10642__A2 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05849__I _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09260__A2 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11323_ _05162_ _05163_ _05164_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11254_ _05000_ _05004_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10704__B _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ _03952_ _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11185_ _04856_ _04923_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10136_ net103 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10067_ _03797_ _03800_ _03802_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_47_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08523__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08523__B2 _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10330__A1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09079__A2 _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10969_ _04707_ _04710_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06837__A1 _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05759__I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06160_ _05348_ _05372_ _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06091_ _05301_ _05305_ _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09850_ _03483_ _03543_ _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07565__A2 _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08801_ _02284_ _02426_ _02427_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09781_ _03407_ _03490_ _03491_ _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06993_ _00470_ _00497_ _00519_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08732_ _02351_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05944_ _03988_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08663_ _02274_ _02275_ _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_94_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05875_ _03226_ _03237_ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ _01135_ _01136_ _01137_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input119_I b_operand[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08594_ _00790_ _00815_ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07545_ _00843_ _01040_ _01064_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_50_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07476_ _00996_ _00997_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_22_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__A2 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06427_ _05561_ _05636_ _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09215_ _02853_ _02875_ _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ _02798_ _02800_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input84_I b_operand[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06358_ _05329_ _05565_ _05568_ _05569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08045__A3 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09077_ _02653_ _02660_ _02664_ _02667_ _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_135_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09793__A3 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06289_ _05499_ _05500_ _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08028_ _01584_ _01586_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07556__A2 _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09979_ _03706_ _03707_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_39_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10823_ _04363_ _04620_ _04621_ _04511_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_72_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08808__A2 _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10754_ _04545_ _04546_ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09481__A2 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10685_ _04400_ _00049_ _05591_ _04472_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07794__I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08992__A1 _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11306_ _05088_ _05108_ _05145_ _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11237_ _05069_ _05070_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08744__A1 _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11168_ net104 _04257_ _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10119_ net106 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11099_ _04869_ _04921_ _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07330_ _00852_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10609__B _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ net72 _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09000_ _02638_ _02641_ _02642_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06212_ _04107_ _05318_ _05355_ _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07192_ _00715_ _00716_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09224__A2 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06143_ _05355_ _05356_ _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06038__A2 _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07235__A1 _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06074_ _05288_ _03171_ _04702_ _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09902_ _03287_ _02333_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07538__A2 _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07209__I _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09833_ _03362_ _03434_ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06113__I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07943__C1 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06210__A2 _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09764_ _03376_ _03431_ _03472_ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06976_ _00502_ _00503_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05952__I _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08715_ _02332_ _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05927_ _02346_ _03759_ _03781_ _03803_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09695_ _03395_ _03397_ _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05858_ _02932_ _02986_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08646_ _02256_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08577_ _00933_ _00872_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05789_ net88 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07528_ _00736_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09463__A2 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07474__A1 _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07459_ _00957_ _00962_ _00861_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10470_ _04198_ _04230_ _04239_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_output190_I net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09129_ _02782_ _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07777__A2 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10781__A1 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11022_ _04834_ _04837_ _01488_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10533__A1 _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06201__A2 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11089__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07701__A2 _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10806_ _04234_ _03912_ _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07465__A1 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06268__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10737_ _04380_ _04526_ _04527_ _04445_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__07465__B2 _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10668_ _04369_ _04372_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11013__A2 _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10599_ _04195_ _03939_ _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10524__A1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09390__A1 _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06830_ _00271_ _00282_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06868__I _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05772__I _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07940__A2 _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06761_ net24 net78 _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09142__A1 _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08500_ _02094_ _02099_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05712_ _01433_ _01444_ _01455_ _01466_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__10827__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09480_ _03096_ _03109_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06692_ _02118_ _03824_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08431_ _01954_ _01959_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08362_ _01935_ _01949_ _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07313_ _00835_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08293_ _01867_ _01874_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07244_ _00766_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07471__A4 _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07208__A1 _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07175_ _00648_ _00660_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06126_ _03171_ _05286_ _03335_ _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06057_ _05213_ _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input47_I a_operand[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10515__A1 _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09381__A1 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09381__B2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ _03423_ _03425_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05682__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09747_ _02556_ _03452_ _03454_ _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06959_ _00373_ _00378_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09133__A1 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10818__A2 _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08993__I _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09678_ _03303_ _03332_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09684__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A1 _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output203_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08629_ _02239_ _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__A1 _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10046__A3 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07447__B2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10451__B1 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10522_ _03904_ _04295_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10453_ _00137_ _04173_ _04208_ _02812_ _04221_ net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_108_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__A1 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10384_ _03976_ _05180_ _04145_ _04146_ _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08175__A2 _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11005_ _04817_ _04637_ _02692_ _04819_ _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10809__A2 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09675__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07686__A1 _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09427__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07312__I _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07438__A1 _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11234__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07989__A2 _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06661__A2 _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05767__I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08938__A1 _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08980_ _02581_ _00049_ _01368_ _02613_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07931_ _01353_ _01327_ _01481_ _01403_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_111_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09363__A1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06177__A1 _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07862_ _01341_ _01331_ _01347_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_68_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11170__A1 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11170__B2 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09601_ _03105_ _03293_ _03294_ _03295_ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_06813_ _00296_ _00299_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07793_ _00979_ _01331_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09532_ _03044_ _03220_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06744_ _00110_ _00273_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09463_ _02458_ _03053_ _00989_ _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06675_ _02291_ _02335_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input101_I b_operand[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08414_ _02002_ _02005_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09394_ _02642_ _03069_ _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09418__A2 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07222__I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07429__A1 _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08345_ _01930_ _01931_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07429__B2 _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08276_ _05431_ _01856_ _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07227_ _00750_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06652__A2 _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08929__A1 _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05677__I _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07158_ _00604_ _00663_ _00682_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10736__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10736__B2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06109_ _03269_ _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06404__A2 _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07601__A1 _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07089_ _02140_ _05365_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08988__I _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output153_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09354__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07904__A2 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09106__A1 _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__B2 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10758__I _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__B1 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10975__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10493__I _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10505_ _04030_ _04276_ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07840__A1 _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06643__A2 _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07840__B2 _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10436_ _04199_ _04202_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08396__A2 _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10367_ _03976_ _05191_ _05267_ _04066_ _04128_ _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10298_ _03823_ _04055_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09345__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11152__A1 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07307__I _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09648__A2 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07659__A1 _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08320__A2 _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06460_ _05609_ _05667_ _05668_ _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06391_ _05596_ _05600_ _05601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06882__A2 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08130_ _01610_ _01614_ _01697_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08084__A1 _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08061_ _00738_ _00786_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07012_ _02401_ _02532_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08387__A2 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06398__A1 _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08963_ _02517_ _02562_ _02566_ _02569_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_25_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09336__A1 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07914_ _01457_ _01460_ _01462_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09336__B2 _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08894_ _02525_ _02528_ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07898__A1 _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07845_ _01378_ _01387_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10497__A3 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ _01163_ _01311_ _01312_ _01231_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_25_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05960__I _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09515_ _03188_ _03201_ _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06727_ _03683_ _02802_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09446_ _03122_ _03123_ _03126_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06658_ _00161_ _00187_ _00188_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06322__A1 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09377_ _02459_ _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06589_ _00119_ _00120_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08328_ _01838_ _01843_ _01913_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08259_ _01718_ _00845_ _00750_ _00785_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11270_ _05089_ _05107_ _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10221_ _03952_ _03960_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10152_ _03894_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10083_ _03819_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11134__A1 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09878__A2 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07889__A1 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10488__A3 _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05870__I _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10985_ _04794_ _04797_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06187__B _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08302__A2 _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06313__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07797__I _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08066__A1 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10948__A1 _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09802__A2 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10419_ _04112_ _04184_ _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11399_ _05155_ _05247_ _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10176__A2 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05960_ _04161_ _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11125__A1 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09869__A2 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05891_ _03378_ _03411_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_94_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08541__A2 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07630_ _01101_ _01105_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05780__I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07561_ _01024_ _01062_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_34_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09300_ _02297_ _01251_ _02960_ _01255_ _02968_ _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_94_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06512_ _01412_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ _00851_ _00763_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06304__A1 _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06304__B2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09231_ _01152_ _02882_ _02885_ _02580_ _02893_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06443_ _05652_ _05653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09162_ _02818_ _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06374_ _05519_ _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08113_ _01675_ _01678_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09093_ _01727_ _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08044_ _01523_ _01527_ _01603_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09557__A1 _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11364__A1 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09995_ _02282_ _02624_ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _02584_ _00240_ _02396_ _01035_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06791__A1 _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08877_ _02490_ _02491_ _02509_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_29_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07828_ _01300_ _01367_ _01369_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_45_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05690__I _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07759_ _01221_ _01225_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08296__A1 _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10770_ _04108_ _04562_ _04563_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__A3 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09429_ _03100_ _03108_ _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07410__I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11322_ _03859_ _03904_ _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09548__A1 _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11253_ _04965_ _04977_ _04975_ _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10204_ _03951_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11184_ _04858_ _04922_ _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10135_ _03870_ _03873_ _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09781__B _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08771__A2 _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10066_ _03699_ _03720_ _03801_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08523__A2 _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09720__A1 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10881__A3 _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10968_ _04704_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08826__A3 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06837__A2 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10899_ _03898_ _04433_ _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07320__I _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10397__A2 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06090_ _05136_ _05303_ _05304_ _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _02278_ _02283_ _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09780_ _02245_ _02431_ _03423_ _03410_ _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06992_ _00475_ _00496_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _02350_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05943_ _02096_ _03955_ _03977_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08662_ net62 _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_54_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06525__A1 _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05874_ net81 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07613_ _00942_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08593_ _00921_ _00905_ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07544_ _00985_ _00981_ _00841_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08278__A1 _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07475_ _00953_ _00847_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09214_ _02863_ _02874_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06426_ _05559_ _05563_ _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07230__I _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09145_ _02795_ _02799_ _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06357_ _05360_ _05223_ _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08986__C1 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input77_I b_operand[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09076_ _02720_ _02724_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06288_ _05440_ _05432_ _05449_ _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08027_ _01579_ _00787_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05685__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07005__A2 _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09950__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09978_ _02462_ _02359_ _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06764__A1 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08929_ _02374_ _02249_ _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08505__A2 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07405__I _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10822_ _03879_ _03958_ _03811_ _03868_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09466__B1 _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10753_ _04413_ _04462_ _04460_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06819__A2 _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10684_ _04471_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08441__A1 _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11305_ _05056_ _05087_ _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08992__A2 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11236_ _04614_ _04214_ _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08744__A2 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11167_ _04980_ _04994_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06755__A1 _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10118_ _03853_ _03857_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11098_ _04873_ _04920_ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10049_ _03238_ _02342_ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07315__I _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07180__A1 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07260_ _00782_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06211_ _05420_ _05421_ _05423_ _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_07191_ _00619_ _00625_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06142_ _04822_ _02672_ _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07235__A2 _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10625__B _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06073_ _02878_ _03117_ _05288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11319__A1 _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06994__A1 _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09901_ _02891_ _03622_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09832_ _03365_ _03432_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06746__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07943__B1 _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06746__B2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07943__C2 _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09763_ _03379_ _03380_ _03430_ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06975_ _00429_ _00430_ _00501_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input131_I b_operand[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08714_ _02331_ _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05926_ _02194_ _03792_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09694_ _02818_ _03393_ _03396_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07225__I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08645_ _02255_ net128 _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05857_ _01260_ _01281_ _02031_ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10845__A3 _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08576_ _00778_ _00822_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05788_ _02291_ _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10058__A1 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07527_ _01045_ _01046_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08120__B1 _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__A3 _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07458_ _00957_ _00972_ _00962_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_50_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11007__B1 _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06409_ _05564_ _05570_ _05618_ _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07389_ _00911_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09128_ net119 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output183_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08423__A1 _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09059_ _02559_ _02592_ _02648_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11021_ _04016_ _04108_ _04836_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06737__A1 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10533__A2 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09687__B1 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10049__A1 _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10805_ _03907_ _04214_ _04446_ _04235_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10736_ _03908_ _03926_ _03939_ _04237_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07465__A2 _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10667_ _03943_ _03873_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08414__A1 _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10598_ _04232_ _04376_ _04378_ _04308_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10221__A1 _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09914__A1 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11219_ _05048_ _05051_ _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10524__A2 _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06760_ _02172_ _01998_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05951__A2 _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05711_ _01184_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10288__A1 _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06691_ _00138_ _00146_ _00221_ net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08430_ _01920_ _01932_ _01930_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08361_ _01943_ _01948_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07312_ _00834_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08292_ _01873_ _01769_ _00937_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10460__A1 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07243_ _00765_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07208__A2 _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07174_ _00642_ _00661_ _00698_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06125_ _05288_ _05286_ _05338_ _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06056_ net15 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06719__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05963__I _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09815_ _03314_ _03527_ _03528_ _03408_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09381__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ _03453_ _02829_ _02555_ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06958_ _02401_ net19 _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05942__A2 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09133__A2 _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05909_ _02456_ _02521_ _03607_ _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ _03377_ _03331_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06889_ _02085_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08628_ _02230_ _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A2 _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08559_ _02109_ _02113_ _02163_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__A2 _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10521_ _03840_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10451__A1 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10451__B2 _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10452_ _03910_ _02744_ _04211_ _04213_ _04220_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_109_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08947__A2 _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10383_ _03975_ _05583_ _04143_ _02692_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10754__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05873__I _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11004_ _04818_ _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08883__A1 _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05697__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07438__A2 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10719_ _03818_ _03866_ _03877_ _03811_ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06949__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10745__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06413__A3 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07610__A2 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07930_ _01402_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05783__I _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07861_ _05104_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07374__A1 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09600_ _02333_ _03014_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06812_ _00296_ _00299_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07792_ _01253_ _01261_ _01272_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09531_ _03135_ _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06743_ _02401_ net17 _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09462_ _02964_ _00235_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06674_ _00149_ _00204_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08413_ _02003_ _02004_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_91_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09393_ _02466_ _03062_ _03068_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08344_ _01925_ _01929_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07429__A2 _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10433__A1 _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08275_ _01680_ _01688_ _01767_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10984__A2 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05958__I _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07226_ _00749_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08929__A2 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05860__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07157_ _00606_ _00662_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10736__A2 _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06108_ _05318_ _01651_ _03248_ _05320_ _05322_ _05323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07601__A2 _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07088_ _00363_ _00612_ _00613_ _00528_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06039_ _04995_ _05006_ _05017_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_59_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05693__I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10104__I _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07614__S _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A2 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09729_ _03265_ _03336_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__A1 _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__B2 _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A2 _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06029__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09290__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10975__A2 _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10504_ _04168_ _04274_ _04275_ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10435_ _04184_ _04200_ _04201_ _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09042__A1 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10366_ _00395_ _04127_ _03963_ _04366_ _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10297_ _04053_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07356__A1 _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07323__I _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06331__A2 _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06390_ _04713_ _05598_ _05599_ _05600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08084__A2 _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08060_ _00913_ _01089_ _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07011_ _00524_ _00537_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09033__A1 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07595__A1 _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08962_ _02562_ _02600_ _02601_ _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_88_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07913_ _01127_ _01458_ _01461_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09336__A2 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08893_ _02526_ _02527_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07844_ _01383_ _01386_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_57_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07898__A2 _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07775_ _00824_ _00846_ _00751_ _00889_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06570__A2 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09514_ _02793_ net61 _03119_ _02484_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_71_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06726_ _00161_ _00188_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08847__A1 _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07233__I _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ _03124_ _03125_ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06657_ _03683_ net78 _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A2 _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09376_ _01118_ _03050_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06588_ _00063_ _00064_ _00117_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10594__I _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08327_ _01840_ _01911_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10957__A2 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08258_ _01729_ _01834_ _01837_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07209_ _04626_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08189_ _01761_ _01762_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08999__I _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10220_ _03823_ _03844_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08378__A3 _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10543__B _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10151_ _03893_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07408__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10082_ _03818_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07338__A1 _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11134__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10984_ _04793_ _04795_ _04796_ _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_74_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10645__A1 _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07510__A1 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08066__A2 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09015__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10418_ _04183_ _03957_ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11398_ _05160_ _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07577__A1 _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10349_ _04106_ _04108_ _04109_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07041__A3 _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11125__A2 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05890_ _03400_ _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07560_ _00999_ _01019_ _01061_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_65_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06511_ _00043_ _05646_ _05652_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07491_ _00864_ _01010_ _05663_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06304__A2 _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _02888_ _02892_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06442_ _05651_ _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09161_ _02318_ _02322_ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09254__A1 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06373_ _03574_ _02510_ _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08112_ _01676_ _01677_ _00944_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06068__A1 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11061__A1 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09092_ _02740_ _02742_ _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_107_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ _00757_ _01489_ _01528_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08612__I _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09557__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10363__B _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ _03608_ _03630_ _03723_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07228__I _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06240__A1 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08945_ _02394_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06791__A2 _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08876_ _02508_ _02386_ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05971__I _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10324__B1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input22_I a_operand[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07827_ _00737_ _00799_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07758_ _01222_ _01224_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10627__A1 _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06709_ _00210_ _03824_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09493__A1 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ _01160_ _01217_ _01218_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _03103_ _03107_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_40_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__A4 _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09359_ _02665_ _02290_ _02300_ _02938_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09245__A1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11321_ _03989_ _03893_ _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11252_ _05056_ _05087_ _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09548__A2 _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10203_ _03950_ _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11183_ _04937_ _04941_ _05012_ _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_121_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08220__A2 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10134_ _03870_ _03874_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10065_ _03670_ _03697_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10866__A1 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10967_ _04765_ _04777_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09484__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08287__A2 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08826__A4 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10898_ _04673_ _04700_ _04703_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_31_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09236__A1 _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09539__A2 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06470__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06991_ _00515_ _00517_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ net53 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05942_ _03966_ _02085_ _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05791__I _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08661_ _02273_ _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05873_ _03215_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06525__A2 _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07612_ _00869_ _01039_ _00882_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10202__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08592_ _02198_ _02099_ _02199_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07543_ _01024_ _01062_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09475__A1 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08278__A2 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06836__B _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11282__A1 _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07474_ _00993_ _00995_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09213_ _02866_ _02868_ _02873_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_139_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06425_ _04822_ _02379_ _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09144_ _02595_ _02323_ _02340_ _02658_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_06356_ _05414_ _05565_ _05566_ _05480_ _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07789__A1 _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08986__B1 _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09075_ _02616_ _02721_ _02723_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08986__C2 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06287_ _05440_ _05432_ _05449_ _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__09438__I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06461__A1 _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08026_ _00782_ _00787_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11337__A2 _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09950__A2 _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09977_ _02433_ _02348_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08928_ _02388_ _02563_ _02565_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09163__B1 _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09702__A2 _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10848__A1 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10848__B2 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08859_ _02224_ _02475_ _02238_ _02240_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10112__I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10821_ _03866_ _04375_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09466__A1 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09466__B2 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10752_ _04497_ _04544_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10683_ _03869_ _03873_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09218__A1 _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08961__B _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11025__A1 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11025__B2 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08441__A2 _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05876__I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11304_ _05140_ _05143_ _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11328__A2 _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11235_ _04004_ _04446_ _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06204__A1 _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11166_ _04989_ _04993_ _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07952__A1 _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06755__A2 _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10117_ _03855_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11097_ _04892_ _04918_ _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10048_ _02267_ _02624_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07180__A2 _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11264__A1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09209__A1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06210_ _05234_ _04550_ _05366_ _05422_ _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__11016__A1 _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06691__A1 _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07190_ _00614_ _00618_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06141_ _05304_ _05351_ _05354_ _04995_ _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05786__I _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06072_ _05286_ _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09900_ _02298_ _02782_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09831_ _03546_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07943__A1 _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07943__B2 _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09762_ _03374_ _03375_ _03373_ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06974_ _00429_ _00430_ _00501_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08713_ net118 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05925_ _02237_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09693_ _02312_ _02332_ _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input124_I b_operand[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08644_ net64 _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05856_ _03019_ _03030_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07171__A2 _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ _02122_ _02179_ _02180_ _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05787_ _02280_ _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11255__A1 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07526_ _01016_ _01018_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09999__A2 _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07241__I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08120__A1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__B2 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07457_ _01423_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06408_ _05567_ _05569_ _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11007__A1 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11007__B2 _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07388_ net6 _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09127_ _02334_ _02235_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06339_ _05548_ _05549_ _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08423__A2 _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05696__I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10230__A2 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09058_ _02677_ _02682_ _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output176_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08009_ _01530_ _01566_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11020_ _04027_ _04051_ _04835_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07934__A1 _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06737__A2 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07416__I _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09687__B2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07698__B1 _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09151__A3 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10049__A2 _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11246__A1 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10804_ _04587_ _04599_ _04600_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_25_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10735_ _04374_ _04441_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10666_ _04368_ _04383_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10597_ _03909_ _03958_ _03812_ _03899_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06425__A1 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11218_ _04961_ _05050_ _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08710__I _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11149_ _04969_ _04974_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05710_ _01173_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06690_ _05666_ _00205_ _00209_ _05317_ _00220_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08360_ _01945_ _01946_ _01947_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08102__A1 _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07061__I _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07311_ _00833_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08291_ _00932_ _00935_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07242_ _00764_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06664__A1 _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10460__A2 _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07173_ _00697_ _00641_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08405__A2 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09602__A1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06124_ _03226_ _05325_ _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06055_ _01401_ _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__A1 _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08620__I _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07916__A1 _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06719__A2 _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09814_ _03406_ _03409_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_59_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09745_ _02276_ _02440_ _02441_ _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06957_ _00471_ _00484_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05908_ _02629_ _03531_ _03542_ _03596_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09676_ _03307_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06888_ _02063_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08627_ _02236_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05839_ _02845_ _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08892__A2 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08558_ _02105_ _02162_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07509_ _01029_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08489_ _01994_ _01999_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09841__A1 _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10520_ _04230_ _04292_ _04293_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06655__A1 _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10451_ _04388_ _04033_ _04217_ _00959_ _04219_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_108_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10382_ _03915_ _00130_ _00394_ _04080_ _04144_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_136_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06958__A2 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07907__A1 _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11003_ _03853_ _04728_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08332__A1 _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08332__B2 _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08883__A2 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05697__A2 _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06646__A1 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ _03865_ _03810_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08705__I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10649_ _04433_ _03931_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09060__A2 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06949__A2 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _01354_ _01404_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07374__A2 _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06811_ _00337_ _00338_ _00339_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07791_ _01253_ _01261_ _01273_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09530_ _03136_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06742_ _00173_ _00177_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07126__A2 _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09461_ _03141_ _03143_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06673_ _00152_ _00203_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10210__I _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08412_ _01718_ _00819_ _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06885__A1 _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09392_ _02288_ _02293_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08343_ _01925_ _01929_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10433__A2 _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08274_ _01767_ _01680_ _01688_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08615__I _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10366__B _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ net16 _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07156_ _00593_ _00679_ _00680_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09051__A2 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06107_ _03324_ _01227_ _05321_ _05287_ _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07087_ _00525_ _00529_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07062__B2 _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input52_I a_operand[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05974__I _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06038_ _01119_ _02824_ _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09354__A3 _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08562__A1 _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output139_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07989_ _00893_ _01096_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ _03362_ _03434_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_47_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09659_ _03358_ _03339_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__A2 _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10120__I _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09814__A1 _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06628__A1 _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10503_ _03982_ _04168_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10434_ _03940_ _03951_ _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09042__A2 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07053__A1 _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10365_ _03965_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09356__I _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10296_ _04052_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11137__B1 _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07356__A2 _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09305__B _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08856__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08608__A2 _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07010_ _00531_ _00536_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05794__I _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08961_ _02518_ _02561_ _02598_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10205__I _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07912_ _00884_ _00877_ _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08892_ _02475_ _02381_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07843_ _01380_ _01384_ _01385_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_69_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10351__A1 _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07774_ _00894_ _01088_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07514__I _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ _02244_ _02430_ _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06725_ _00185_ _00197_ _00254_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08847__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06858__A1 _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09444_ _02512_ net59 net58 _02249_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06656_ net24 net77 _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06587_ _00065_ _00118_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09375_ _02959_ _02961_ _02466_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05969__I _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08326_ _01262_ _01835_ _01841_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08257_ _01630_ _01835_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07208_ _00678_ _00731_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08188_ _01695_ _01696_ _01759_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07035__A1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07139_ _00593_ _00596_ _00664_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_106_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08783__A1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06389__A3 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _03892_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10590__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10115__I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10081_ net30 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10342__A1 _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10983_ _04393_ _03907_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06849__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07510__A2 _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09263__A2 _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10417_ _03931_ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11397_ _05167_ _05179_ _05244_ _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07577__A2 _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08774__A1 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10348_ _04074_ _04089_ _04053_ _03968_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10279_ _03906_ _04034_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10333__A1 _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06510_ _03672_ _03727_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07490_ _00864_ _01010_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06441_ _02379_ _02434_ _05651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05789__I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09160_ _02316_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06372_ _05279_ _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09254__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08111_ _00788_ _00927_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06068__A2 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09091_ _02646_ _02685_ _02741_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11061__A2 _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08042_ _01516_ _01600_ _01601_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09006__A2 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07017__A1 _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08114__B _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07509__I _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09993_ _03612_ _03628_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08944_ _02581_ _05191_ _05267_ _02402_ _02582_ _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08517__A1 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _02507_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10324__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10324__B2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07826_ _00813_ _01088_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input15_I a_operand[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05751__A1 _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ _00746_ _00804_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10627__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06708_ _01803_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ _01215_ _01166_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09493__A2 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ _03101_ _03104_ _03105_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_80_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06639_ _03640_ _05353_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09358_ _02939_ _02941_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09245__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08309_ _01787_ _01791_ _01892_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07256__A1 _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09289_ _02461_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11320_ _04005_ _03914_ _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08803__I _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11251_ _05075_ _05086_ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08756__A1 _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ _03949_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11182_ _04950_ _05011_ _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _03873_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07863__B _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10064_ _03728_ _03729_ _03799_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10315__A1 _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09181__A1 _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10866__A2 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__A2 _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10966_ _04770_ _04776_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10897_ _04701_ _03948_ _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08713__I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06470__A2 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08747__A1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06233__I _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06990_ _00454_ _00516_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input7_I a_operand[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05941_ _02063_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05981__A1 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08660_ _02272_ _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05872_ _03204_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09711__A3 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07611_ _01041_ _01039_ _01134_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08591_ _02089_ _02093_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07542_ _01020_ _01061_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10609__A2 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07473_ _00956_ _00994_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09212_ _02864_ _02869_ _02870_ _02871_ _02872_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06424_ _05558_ _05571_ _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07238__A1 _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09143_ _02228_ _02325_ _02341_ _02485_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06355_ _02715_ _02921_ _01553_ _03411_ _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08986__A1 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09074_ _02358_ _02722_ _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08986__B2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08623__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06286_ _05497_ _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__A3 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08025_ _01345_ _01507_ _01571_ _01406_ _01583_ net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_144_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07239__I _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09976_ _02267_ _02393_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08927_ _02230_ _02376_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09163__B2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08858_ _02483_ _02490_ _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10848__A2 _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07809_ _00818_ _01348_ _01274_ _00908_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_55_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08789_ _02343_ _02354_ _02411_ _02414_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_72_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10820_ _04613_ _04618_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09466__A2 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10751_ _04500_ _04543_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10682_ _03994_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11025__A2 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08977__A1 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11303_ _05141_ _05142_ _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06452__A2 _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11234_ _03987_ _03903_ _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06053__I _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10536__A1 _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06204__A2 _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07401__A1 _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11165_ _04990_ _04991_ _04992_ _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_1_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05892__I _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07952__A2 _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10116_ _03854_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11096_ _04893_ _04917_ _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_48_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10047_ _03622_ _03758_ _03714_ _03712_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10303__I _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10839__A2 _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08901__A1 _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07468__A1 _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10949_ _04685_ _04758_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07468__B2 _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09209__A2 _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06140_ _02813_ _05353_ _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08968__A1 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06071_ _03291_ _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10922__B _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09393__A1 _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09830_ _03471_ _03545_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07943__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09761_ _03464_ _03469_ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06973_ _00432_ _00435_ _00500_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09145__A1 _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ _02321_ _02329_ _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05924_ _03770_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09692_ _03181_ _03393_ _03394_ _03297_ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ _02253_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05855_ _02020_ _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input117_I b_operand[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08574_ _02124_ _02137_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08618__I _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09448__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05786_ _02269_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07525_ _00993_ _01017_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07459__A1 _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08120__A2 _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07456_ _00972_ _00976_ _00977_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06138__I _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06407_ _05555_ _05616_ _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11007__A2 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07387_ _00802_ _00808_ _00909_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_input82_I b_operand[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08959__A1 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09126_ _02221_ _02320_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06338_ _05471_ _05474_ _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06074__S _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09057_ _02454_ _02703_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06269_ net82 _05352_ _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _01532_ _01549_ _01565_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_116_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output169_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06198__A1 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09959_ _02277_ _03014_ _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10123__I _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09687__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10803_ _03871_ net96 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05712__A4 _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10734_ _04522_ _04523_ _04524_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__06048__I _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10665_ _04429_ _04432_ _04450_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_40_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05887__I _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10596_ _04374_ _04375_ _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06425__A2 _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08178__A2 _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11217_ _04959_ _04964_ _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09094__I _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07925__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11148_ _04969_ _04974_ _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_110_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05936__A1 _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09127__A1 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11079_ _03987_ _04441_ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11237__A2 _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07310_ net102 _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08290_ _00940_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07241_ net80 _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05797__I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07172_ _00608_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06123_ _05336_ _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06054_ _04312_ _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11173__A1 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09813_ _03114_ _02625_ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09744_ _02441_ _03251_ _02276_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06956_ _00479_ _00483_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_74_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05907_ _03574_ _03585_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09675_ _03374_ _03375_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06887_ _03966_ _00414_ _04269_ _00231_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__A2 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08626_ _02235_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05838_ _02834_ _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06352__A1 _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07252__I _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ _02114_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05769_ _02063_ _02085_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07508_ net38 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08488_ net75 _00844_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07852__A1 _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07439_ _00740_ _00756_ _00769_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06655__A2 _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10450_ _04218_ _00232_ _00131_ _03917_ _04258_ _03976_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__10739__A1 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09109_ _02471_ _02760_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07604__A1 _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11400__A2 _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ _05202_ _04143_ _03929_ _00397_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_108_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09357__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07907__A2 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11002_ _04816_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09109__A1 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08580__A2 _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07135__A3 _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06343__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08883__A3 _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11219__A2 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06894__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08096__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10978__A1 _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10717_ _03818_ _03987_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06646__A2 _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10648_ _04257_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10579_ _04296_ _04300_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09348__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09899__A2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08571__A2 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06810_ _00264_ _00283_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07790_ _01326_ _01328_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06741_ _00265_ _00270_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08859__B1 _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09460_ _05375_ _03142_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06672_ _00154_ _00202_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08411_ _00784_ _00870_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09391_ _02460_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08342_ _01926_ _01928_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10969__A1 _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07834__A1 _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08273_ _01777_ _01853_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10366__C _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07224_ _00745_ _00747_ _01498_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07155_ _00594_ _00595_ _00664_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06106_ _01357_ _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07086_ _02074_ _02889_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07062__A2 _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06037_ _02921_ _02009_ _05006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11146__A1 _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07247__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input45_I a_operand[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06151__I _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08562__A2 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07988_ _00809_ _00874_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06573__A1 _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09727_ _03365_ _03432_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06939_ _00461_ _00465_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09658_ _03156_ _03217_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08609_ _02152_ _02217_ _02218_ _00735_ net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_output201_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09589_ _03180_ _03183_ _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08078__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08806__I _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06527__S _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07825__A1 _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _03981_ _04267_ _03906_ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10433_ _03926_ _03841_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10364_ _03967_ _04125_ _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11137__A1 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10295_ _04027_ _04051_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11137__B2 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08002__A1 _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09750__A1 _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07513__B1 _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08716__I _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09569__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08241__A1 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08960_ _02230_ _02364_ _02388_ _02568_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_88_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07911_ _01315_ _01458_ _01459_ _01384_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_102_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08891_ _02245_ _02239_ _02254_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08544__A2 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__A1 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07842_ net124 _01074_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09741__B2 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07773_ _01306_ _01309_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09512_ _03194_ _03198_ _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06724_ _00186_ _00196_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09443_ _02595_ _03120_ _02299_ _02484_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_92_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06655_ _00108_ _00111_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09374_ _03048_ _02959_ _02961_ _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08626__I _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06586_ _00117_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07530__I _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08325_ _01809_ _01817_ _01909_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07807__A1 _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08256_ _00797_ _01156_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06146__I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07207_ _00678_ _00731_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08187_ _01695_ _01696_ _01759_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11367__A1 _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08232__A1 _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07138_ _00604_ _00663_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07035__A2 _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07069_ _00518_ _00570_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06794__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10590__A2 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output151_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10080_ _03816_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10840__B _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09732__A1 _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06546__A1 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08299__A1 _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10982_ net40 net98 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06849__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09799__A1 _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06056__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10416_ _04124_ _04155_ _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11396_ _05153_ _05166_ _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10030__A1 _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08774__A2 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10347_ _04052_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06785__A1 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10278_ _03981_ _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08526__A2 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07615__I _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06440_ _03705_ _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07350__I _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06371_ _05580_ _05581_ _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08110_ _01588_ _01589_ _00788_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07265__A2 _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09090_ _02573_ _02609_ _02684_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08041_ _01519_ _01568_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11349__A1 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06225__B1 _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09992_ _03667_ _03721_ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10572__A2 _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08943_ _00395_ _02396_ _02395_ _00397_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08517__A2 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09714__A1 _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08874_ _02225_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06528__A1 _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07725__B1 _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10324__A2 _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07825_ _01302_ _01319_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ _01214_ _01289_ _01290_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05751__A2 _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06707_ _05319_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07687_ _01215_ _01166_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09426_ _02318_ _02625_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06638_ _00101_ _00104_ _00112_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07260__I _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06700__A1 _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09357_ _03027_ _03029_ _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06569_ _03661_ _03019_ _00100_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ _00756_ _00931_ _01793_ _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__A2 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09288_ _02897_ _02955_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output199_I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08239_ _01812_ _01816_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11250_ _05078_ _05085_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07008__A2 _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10201_ _03948_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09953__A1 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11181_ _04953_ _05010_ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06767__A1 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10132_ _03872_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09705__A1 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10063_ _03798_ _03726_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06519__A1 _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09181__A2 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10965_ _04772_ _04775_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10896_ net41 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08444__A1 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08747__A2 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11379_ _05170_ _05178_ _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05940_ _03845_ _03922_ _03944_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05871_ _03193_ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09711__A4 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07183__A1 _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07610_ _00873_ _01072_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08590_ _02094_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07541_ _01047_ _01060_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07472_ _00738_ _00851_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09211_ _02864_ _02869_ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06423_ _05617_ _05619_ _05632_ _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_22_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09142_ _02792_ _02796_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08435__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08904__I _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07238__A2 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06354_ _05477_ _02899_ _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09073_ _02514_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08986__A2 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06285_ _01727_ _05497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08024_ _01500_ _05644_ _01574_ _05648_ _01582_ _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_89_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06749__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10545__A2 _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09975_ _03594_ _03602_ _03702_ _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08926_ _02250_ _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09163__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08857_ _02488_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07808_ _01269_ _01271_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08910__A2 _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08788_ _02337_ _02413_ _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06921__A1 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07739_ _01272_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10750_ _04503_ _04542_ _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09409_ _02746_ _03015_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06685__B1 _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10681_ _04467_ _04468_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_138_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08977__A2 _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08035__B _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06988__A1 _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10784__A2 _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11302_ _05094_ _05096_ _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11233_ _05062_ _05066_ _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10536__A2 _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11164_ _04614_ _04446_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07401__A2 _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10115_ net44 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11095_ _04906_ _04916_ _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10046_ _03775_ _03778_ _03779_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_76_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06912__A1 _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10948_ _04688_ _04693_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07468__A2 _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10879_ net105 _04375_ _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06140__A2 _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08417__A1 _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09614__B1 _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10224__A1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06070_ _04930_ _04984_ _05093_ _05115_ _05285_ net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__09917__A1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06600__B1 _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09760_ _03466_ _03468_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06972_ _00444_ _00499_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08711_ _02328_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05923_ _02302_ _02324_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09691_ _02783_ _02340_ _02657_ _03006_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08642_ _02252_ _02235_ _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05854_ _01564_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08573_ _02124_ _02137_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05785_ net24 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07524_ _01040_ _01042_ _05663_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07459__A2 _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10463__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07455_ _00972_ _00976_ _05291_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06406_ _05554_ _05614_ _05615_ _05616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_10_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08408__A1 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08634__I _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07386_ _00818_ _00901_ _00902_ _00908_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10215__A1 _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09125_ _02720_ _02724_ _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06337_ _05472_ _05473_ _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09081__A1 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input75_I b_operand[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09056_ _02354_ _02411_ _02699_ _02702_ _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_68_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06268_ net81 net15 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08007_ _01556_ _01563_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09908__A1 _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06199_ _02694_ _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10518__A2 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07934__A3 _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09958_ _03680_ _03684_ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08909_ _01192_ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07147__A1 _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09889_ _03536_ _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07698__A2 _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08809__I _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06370__A2 _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10802_ net41 net95 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10733_ _03882_ _03949_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10664_ _04437_ _04449_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05881__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09072__A1 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10595_ _03956_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06064__I _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11216_ _04955_ _05046_ _05047_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09375__A2 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11147_ _04970_ _04972_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05936__A2 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09127__A2 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11078_ _04895_ _04896_ _04899_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10029_ _03760_ _03761_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08719__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10445__A1 _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07240_ _00752_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07171_ _00692_ _00695_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09063__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10748__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06122_ _02737_ _03313_ _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06053_ _05169_ _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06702__I _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11173__A2 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ _03514_ _03525_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06955_ _00480_ _00481_ _00482_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09743_ _03441_ _03443_ _03450_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05906_ net85 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09674_ _02435_ _02505_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08877__A1 _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08629__I _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06886_ _05384_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ _02234_ _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05837_ _02824_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08556_ _02078_ _02141_ _02159_ _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05768_ _02074_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07507_ _04086_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08487_ _02083_ _02000_ _02084_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05699_ net3 _01151_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07438_ _00865_ _00950_ _00960_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07369_ net65 _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09108_ _02414_ _02701_ _02343_ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output181_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10380_ _03921_ _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09039_ _02646_ _02685_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07368__A1 _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11164__A2 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11001_ _04020_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06040__A1 _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08868__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07443__I _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06343__A2 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06059__I _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09293__A1 _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08096__A2 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05898__I _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10716_ _04429_ _04504_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10647_ _04373_ _04382_ _04430_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10578_ _04298_ _04299_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07359__A1 _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10902__A2 _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06740_ _00266_ _00267_ _00269_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08859__A1 _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08859__B2 _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09520__A2 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06671_ _00156_ _00201_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07531__A1 _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08410_ _00914_ _00885_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09390_ _02977_ _03047_ _03059_ _03066_ net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_24_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08341_ _01922_ _01927_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08272_ _01779_ _01852_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07834__A2 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07223_ _00740_ _00746_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07154_ _00594_ _00595_ _00664_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07598__A1 _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06105_ _05319_ _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07085_ _00609_ _00530_ _00610_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06270__A1 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06036_ _02965_ _01564_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09339__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input38_I a_operand[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07987_ _01461_ _01540_ _01541_ _01385_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_75_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07770__A1 _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06573__A2 _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09726_ _03376_ _03431_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06938_ _00461_ _00465_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10657__A1 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09657_ _03218_ _03339_ _03340_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_06869_ _00395_ _00396_ _03911_ _00397_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_43_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08608_ _02155_ _02215_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09588_ _03180_ _03183_ _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _02066_ _02069_ _02142_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08078__A2 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09275__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06089__A1 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06607__I _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10501_ _02977_ _04252_ _04264_ _04273_ net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_7_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10129__I _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09027__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10432_ _04196_ _04197_ _04198_ _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ _03971_ _04077_ _04124_ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08250__A2 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06261__A1 _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10294_ _04038_ _04045_ _04050_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__11137__A2 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07882__B _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06013__A1 _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09750__A2 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07513__A1 _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07513__B2 _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__A2 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09266__A1 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11073__A1 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07816__A2 _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10820__A1 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09018__A1 _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08732__I _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07348__I _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07910_ _01380_ _01385_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07792__B _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08890_ _02524_ _02402_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09563__I _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06004__A1 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07841_ _01156_ net113 _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__A2 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07752__A1 _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07772_ _01307_ _01308_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09511_ _03195_ _03196_ _03197_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_37_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06723_ _04107_ _02107_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _02665_ _02279_ _02290_ _02485_ _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06654_ _00090_ _00183_ _00184_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09373_ _02466_ _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06585_ _00068_ _00072_ _00116_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09257__A1 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08324_ _01812_ _01816_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07807__A2 _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ _01723_ _01730_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09009__A1 _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07206_ _00681_ _00683_ _00730_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08186_ _01698_ _01758_ _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11367__A2 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07137_ _00606_ _00662_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07258__I _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07068_ _00520_ _00569_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06794__A2 _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06019_ _01260_ _02997_ _04778_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10878__A1 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08535__A3 _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output144_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07743__A1 _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09709_ _03201_ _03326_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10981_ _04708_ _04792_ _04793_ _04607_ _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_62_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09496__A1 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08299__A2 _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08817__I _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11243__I _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09799__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10802__A1 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06482__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11358__A2 _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08759__B1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10415_ _04158_ _04163_ _04179_ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11395_ _05140_ _05143_ _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10346_ _03954_ _03960_ _04105_ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10030__A2 _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10277_ _03918_ _03974_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09723__A2 _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06537__A2 _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07734__A1 _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07734__B2 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09487__A1 _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08727__I _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07631__I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11046__A1 _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06370_ _05500_ _05514_ _05527_ _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08040_ _01519_ _01568_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09558__I _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06473__A1 _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11349__A2 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08214__A2 _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06225__A1 _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09991_ _03699_ _03720_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08942_ _02364_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07806__I _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09714__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06710__I _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08873_ _02223_ _02505_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07725__A1 _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07824_ _01297_ _01363_ _01364_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07755_ _01220_ _01236_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06706_ _00231_ _00233_ _00234_ _02129_ _00235_ _00129_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_07686_ _01051_ _01163_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08637__I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09425_ net118 net53 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06637_ _00099_ _00166_ _00167_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11037__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09356_ _03028_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06568_ _05359_ _02313_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08307_ _01782_ _01851_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ _02952_ _02953_ _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06499_ _00027_ _00028_ _00031_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08453__A2 _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09650__A1 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06464__A1 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08238_ _01810_ _01813_ _01815_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08169_ _01627_ _01739_ _01740_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10200_ net96 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11180_ _04979_ _05009_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06767__A2 _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ _03871_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09166__B1 _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09705__A2 _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ _03724_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06519__A2 _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10142__I _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09181__A3 _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09469__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10964_ _04768_ _04773_ _04774_ _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_55_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08141__A1 _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10895_ net42 net95 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08444__A2 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11200__A1 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11378_ _05221_ _05204_ _05224_ _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07955__A1 _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10329_ _04060_ _03946_ _04088_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07707__A1 _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05870_ _03182_ _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06930__A2 _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07540_ _01055_ _01059_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07361__I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _00739_ _00851_ _00763_ _00767_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_62_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06422_ _05623_ _05631_ _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09210_ _02326_ _02251_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10490__A2 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09141_ _02795_ _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06353_ _05559_ _05563_ _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09632__A1 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09072_ _02345_ _02486_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06284_ _05104_ _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06705__I _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08023_ _01576_ _01578_ _01580_ _01581_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_135_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10227__I _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08199__A1 _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06749__A2 _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09974_ _03597_ _03601_ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06440__I _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08925_ _02479_ _02516_ _02561_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_58_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09699__A1 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08856_ _02485_ _02487_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_57_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input20_I a_operand[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08371__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07807_ _01337_ _00800_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08787_ _02342_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05999_ _01346_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06382__B1 _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11258__A1 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07738_ _01269_ _01271_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07271__I _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08123__A1 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07669_ _01152_ _01183_ _01185_ _01187_ _01197_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09408_ _02338_ _02344_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06685__A1 _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06685__B2 _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10680_ _04395_ _04391_ _04044_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09339_ _02318_ _02614_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10233__A2 _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11301_ _04960_ _05095_ _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10137__I _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11232_ _05063_ _05065_ _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10536__A3 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11163_ net105 net35 _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10114_ _03852_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11094_ _04910_ _04915_ _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_1_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10045_ _02389_ _03673_ _03674_ _03679_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_64_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08277__I _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10947_ _04695_ _04714_ _04755_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07873__B1 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10878_ _04613_ _04618_ _04627_ _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10756__B _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08417__A2 _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07640__A3 _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09378__B1 _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08740__I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09917__A2 _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06600__A1 _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06971_ _00446_ _00498_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08710_ _02327_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05922_ _02445_ _03618_ _03738_ _03748_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_09690_ _02890_ _02338_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08353__A1 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08641_ _02251_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05853_ _02932_ _02997_ _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06903__A2 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08572_ _02117_ _02138_ _02177_ _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05784_ _02205_ _02247_ _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07523_ _01040_ _01042_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_81_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07454_ _00973_ _00974_ _00975_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10463__A2 _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06405_ _01097_ _02412_ _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07385_ _00905_ _00907_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06419__A1 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11412__A1 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10215__A2 _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06336_ _01303_ _02467_ _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09124_ _02727_ _02775_ _02776_ _02733_ _02725_ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__08959__A3 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09081__A2 _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09055_ _02642_ _02701_ _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06267_ _05361_ _05476_ _05478_ _05415_ _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08006_ _01559_ _01562_ _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input68_I a_operand[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06198_ _05234_ _05409_ _05410_ _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_89_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10923__B1 _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07266__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09957_ _03681_ _03682_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08908_ _02389_ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09888_ _03529_ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08839_ _02455_ _02465_ _02469_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10801_ _04510_ _04514_ _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06107__B1 _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10732_ _03871_ _03840_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ _04444_ _04448_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11403__A1 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07607__B1 _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10594_ _03897_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09072__A2 _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08280__B1 _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11215_ _04958_ _04978_ _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_122_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11146_ _04967_ _04971_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10390__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11077_ _04760_ _04897_ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09391__I _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ _03709_ _03717_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06649__A1 _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08735__I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ _05652_ _00693_ _00694_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09063__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06121_ _05290_ _05293_ _05335_ net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10748__A3 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07074__A1 _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06052_ _01216_ _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06821__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07377__A2 _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09811_ _03519_ _03524_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10381__A1 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09742_ _03351_ _00966_ _03447_ _03449_ _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06954_ _00268_ _05327_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08326__A1 _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07129__A2 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05905_ _03564_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09673_ _03372_ _03373_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08877__A2 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06885_ _05528_ _00409_ _00410_ _00412_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input122_I b_operand[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10240__I _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08624_ _02233_ _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05836_ _02813_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08555_ _02080_ _02139_ _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05767_ net93 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07506_ _00864_ _01026_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08486_ _02001_ _02006_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05698_ net2 _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07437_ _00951_ _00952_ _00958_ _00959_ _00957_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_22_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07368_ _00887_ _00890_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_108_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10739__A3 _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09107_ _01345_ _02705_ _02743_ _01406_ _02758_ net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__07065__A1 _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06319_ _02629_ _03531_ _04951_ _03542_ _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07299_ _00821_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09038_ _02647_ _02684_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_output174_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07368__A2 _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11000_ _04812_ _04814_ _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_120_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08317__A1 _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06591__A3 _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10124__A1 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10150__I _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06879__A1 _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09817__A1 _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09293__A2 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10715_ _04432_ _04450_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07843__A3 _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10646_ _04379_ _04381_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10577_ _03826_ _03883_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07359__A2 _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11129_ _04885_ _04889_ _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08308__A1 _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06582__A3 _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06670_ _00165_ _00200_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_92_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07531__A2 _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09808__A1 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10418__A2 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08340_ _00918_ _00823_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ _01782_ _01851_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07295__A1 _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11091__A2 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07222_ net69 _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09036__A2 _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07153_ _00592_ _00669_ _00677_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08795__A1 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06104_ _01683_ _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07084_ _00531_ _00536_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06035_ _03106_ _04973_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_87_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08011__A3 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07986_ _00888_ _01157_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07770__A2 _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09725_ _03381_ _03430_ _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06937_ _00462_ _00464_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10657__A2 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09656_ _03256_ _03355_ net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06868_ _04366_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08607_ _02155_ _02215_ _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05819_ net18 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09587_ _03277_ _03278_ _03279_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06799_ _00289_ _00300_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05999__I _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ _02078_ _02141_ _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06089__A2 _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08469_ _01983_ _01985_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10500_ _04253_ _04270_ _04272_ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _03820_ _03909_ _03924_ _03812_ _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10362_ _04123_ _03958_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06261__A2 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ _03850_ _04046_ _04047_ _04049_ _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06013__A2 _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07761__A2 _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07513__A2 _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09266__A2 _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09018__A2 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07029__A1 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10629_ _04346_ _04387_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10584__A1 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06252__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08529__A1 _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06004__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07840_ _01232_ _01380_ _01382_ _00878_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_111_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07364__I _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07771_ _00820_ _00834_ _00848_ _00885_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09510_ _02286_ _02385_ _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06722_ _00165_ _00200_ _00251_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09441_ _03028_ _03121_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06653_ _00093_ _00096_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09372_ _02982_ _03046_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06708__I _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06584_ _00081_ _00115_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09257__A2 _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _01819_ _01846_ _01907_ _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08254_ _01821_ _01827_ _01832_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_20_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07205_ _00691_ _00729_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08185_ _01700_ _01757_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06228__C1 _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07136_ _00642_ _00661_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06443__I _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07440__A1 _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07067_ _00515_ _00517_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input50_I a_operand[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06018_ _04778_ _04789_ _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07991__A2 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10590__A4 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09193__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07274__I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07969_ _01451_ _01464_ _01522_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output137_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09708_ _03407_ _03412_ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10980_ _04329_ _04234_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09496__A2 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09639_ _03261_ _03337_ _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10802__A2 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06482__A2 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08759__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10414_ _03943_ _03928_ _04160_ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08759__B2 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11394_ _05189_ _05241_ _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10345_ _03947_ _03962_ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07982__A2 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10276_ _03930_ _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05993__A1 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09184__A1 _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09723__A3 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07734__A2 _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08931__A1 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09487__A2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07498__A1 _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08743__I _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06473__A2 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06225__A2 _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09990_ _03701_ _03719_ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08941_ _05502_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10309__A1 _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09175__A1 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08872_ _02504_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07725__A2 _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07823_ _01291_ _01320_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07754_ _01219_ _01235_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07489__A1 _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06705_ _04258_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07685_ _01049_ _00814_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09424_ _02929_ _03101_ _03102_ _03010_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06636_ _00083_ _00113_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06438__I _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _02225_ _02289_ _02299_ _02476_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_40_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11037__A2 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06567_ _00086_ _00098_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08306_ _01784_ _01850_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input98_I b_operand[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08653__I _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09286_ _02898_ _02900_ _02951_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_60_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06498_ _05621_ _00029_ _00030_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09650__A2 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08237_ _01333_ _01096_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07269__I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08168_ _01554_ _01631_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07119_ _00643_ _00644_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08099_ _01663_ _01664_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10130_ net40 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07964__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10061_ _03774_ _03786_ _03796_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09166__B2 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08913__A1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10720__A1 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08828__I _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10963_ _04512_ _04214_ _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06152__A1 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10894_ _04622_ _04625_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10787__A1 _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10003__A3 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11377_ _05146_ _05222_ _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10328_ _03839_ _04062_ _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09157__A1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10259_ _04012_ _04009_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07707__A2 _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10711__A1 _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08738__I _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07470_ _01847_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09880__A2 _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06421_ _05626_ _05630_ _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_34_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ _02793_ _02339_ _02350_ _02794_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_06352_ _05561_ _05562_ _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09632__A2 _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06283_ _05458_ _05494_ _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09071_ _02221_ _02334_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08022_ _01490_ _05319_ _05519_ _01502_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09396__A1 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09973_ _03617_ _03627_ _03700_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05957__A1 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10950__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08924_ _02560_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09699__A2 _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08855_ _02486_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10702__A1 _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07806_ _05445_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08786_ _02369_ _02405_ _02408_ _02410_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__06382__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08648__I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07552__I _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05998_ _04571_ _02997_ _04495_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input13_I a_operand[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06382__B2 _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11258__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07737_ _01256_ _00807_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08123__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07668_ _01190_ _01194_ _01196_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09407_ _03004_ _03018_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06619_ _00072_ _00116_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06685__A2 _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07599_ _01118_ _01121_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09338_ _02331_ _02625_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09623__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05800__I _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07634__A1 _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ _02796_ _02865_ _02869_ _02934_ _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_138_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11300_ _05092_ _05137_ _05139_ _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11231_ _05059_ _05064_ _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11194__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11162_ net107 _03937_ _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10941__A1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10113_ _03851_ _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06070__B1 _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11093_ _04912_ _04914_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10044_ _03776_ _03693_ _03777_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07462__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11249__A2 _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10946_ _04613_ _04618_ _04627_ _04694_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_44_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07873__A1 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10877_ _04611_ _04678_ _04679_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07873__B2 _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06428__A2 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09378__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09378__B2 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05939__A1 _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06600__A2 _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06970_ _00470_ _00497_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I a_operand[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05921_ _03629_ _03716_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08353__A2 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09550__A1 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08640_ _02250_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05852_ _02986_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07372__I _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _02176_ _02116_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05783_ _02237_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09302__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08105__A2 _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ _01041_ _00869_ _00974_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07453_ _00867_ _00946_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06404_ _02575_ _05353_ _05614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07384_ _00906_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09123_ _02662_ _02732_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06335_ _05466_ _05544_ _05545_ _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10238__I _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07616__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06419__A2 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11412__A2 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08959__A4 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09081__A3 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09054_ _02408_ _02410_ _02640_ _02700_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06266_ _01086_ _05477_ _05360_ _01531_ _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08005_ _01557_ _01560_ _01561_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_135_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06197_ _03204_ _02954_ _05410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10923__A1 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09956_ _03583_ _03589_ _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08907_ _02542_ _01338_ _02403_ _00238_ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09887_ _03502_ _03505_ _03606_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09541__A1 _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08838_ _02437_ _02468_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10687__B1 _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06355__B2 _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07282__I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08769_ _02392_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10800_ _04525_ _04595_ _04596_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06107__A1 _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10731_ _03892_ _04297_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10662_ _04438_ _04445_ _04447_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07607__A1 _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10148__I _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11403__A2 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07607__B2 _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10593_ _04369_ _04372_ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08280__A1 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08841__I _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08280__B2 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07457__I _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11214_ _04958_ _04978_ _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10914__A1 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09780__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11145_ _04701_ _04194_ _04971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10390__A2 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11076_ net109 net31 _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10611__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10027_ _03711_ _03715_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06346__A1 _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10929_ _04662_ _04719_ _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06120_ _05295_ _05313_ _05316_ _05317_ _05334_ _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08751__I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06051_ _03106_ _05147_ _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06821__A2 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11158__A1 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07367__I _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10007__B _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09810_ _03521_ _03522_ _03523_ _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_87_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08574__A2 _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10381__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09741_ _02264_ _05583_ _03448_ _02546_ _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06953_ net87 _02639_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08326__A2 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10521__I _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05904_ _03553_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09672_ _03368_ _03371_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06337__A1 _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06884_ _05444_ _00411_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08877__A3 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08623_ net48 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05835_ _02802_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input115_I b_operand[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08554_ _02066_ _02156_ _02157_ _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05766_ _02053_ _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07505_ _00985_ _00981_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07837__A1 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ _01996_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05697_ _01130_ _01303_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07436_ _05591_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07367_ _00889_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input80_I b_operand[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09106_ _02336_ _02744_ _02750_ _02751_ _02757_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_108_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08661__I _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06318_ _05434_ _02618_ _05393_ _05396_ _05450_ _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07298_ _00820_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09037_ _02677_ _02682_ _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06249_ _05460_ _05426_ _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11149__A1 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07277__I _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08014__A1 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output167_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__A1 _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09939_ _03633_ _03642_ _03663_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09514__A1 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11321__A1 _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10124__A2 _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07828__A1 _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10714_ _04501_ _04457_ _04502_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10645_ _04364_ _04428_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11388__A1 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10576_ _04289_ _04352_ _04353_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_127_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09753__A1 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06567__A1 _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11128_ _04892_ _04918_ _04952_ _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08308__A2 _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11059_ _03854_ _04295_ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09808__A2 _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10823__B1 _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08270_ _01784_ _01850_ _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08492__A1 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07221_ _00742_ _00744_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11379__A1 _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08244__A1 _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07152_ _00665_ _00676_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06103_ _02672_ _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08795__A2 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07598__A3 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07083_ _00527_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06034_ _04940_ _04951_ _04962_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06869__C _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07985_ _01127_ _01458_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_47_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10251__I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09724_ _03402_ _03429_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07770__A3 _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06936_ _00459_ _00463_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_28_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09655_ _03343_ _03347_ _03348_ _03354_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_28_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06867_ _03889_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08606_ _02158_ _02160_ _02214_ _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_43_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05818_ _02564_ _02618_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09586_ _03186_ _03209_ _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08656__I _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06798_ _00289_ _00300_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08537_ _02080_ _02139_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05749_ _01868_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09275__A3 _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08468_ _02062_ _02064_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07419_ _00773_ _00938_ _00941_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08399_ _01935_ _01949_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10430_ _03925_ _03814_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09983__A1 _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10426__I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ _03949_ _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10292_ _04012_ _04048_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06549__A1 _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10805__B1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10281__A1 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10628_ _04346_ _04387_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07029__A2 _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09423__B1 _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10033__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10336__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ _04028_ _05586_ _00133_ _04030_ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06788__A1 _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10584__A2 _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08529__A2 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07770_ _00893_ _01157_ _01087_ _00848_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_49_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05763__A2 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06960__B2 _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06721_ _00168_ _00199_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _02595_ _03119_ _03120_ _02658_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06652_ _00093_ _00096_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07380__I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06712__A1 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09371_ _03044_ _03045_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06583_ _00082_ _00114_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08322_ _01820_ _01845_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08465__A1 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10272__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08253_ _01828_ _01831_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07204_ _00696_ _00699_ _00728_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08184_ _01710_ _01756_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06228__B1 _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10246__I _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__A1 _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07135_ _00646_ _00648_ _00660_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06228__C2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07066_ _00590_ _00591_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07440__A2 _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06017_ _01119_ _04539_ _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09717__A1 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07991__A3 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input43_I a_operand[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09193__A2 _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07968_ _01452_ _01463_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05754__A2 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06951__A1 _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09707_ _03321_ _03410_ _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06919_ _00352_ _00355_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07899_ _01441_ _01445_ _01446_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09638_ _03265_ _03336_ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07290__I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05803__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09569_ _03163_ _03167_ _03260_ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08208__A1 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10413_ _04153_ _04177_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08759__A2 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10156__I _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11393_ _05184_ _05200_ _05240_ _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10344_ _04079_ _04084_ _04104_ net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09708__A1 _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10275_ _04029_ _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10318__A2 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09184__A2 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06942__A1 _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05713__I _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08940_ _02397_ _02578_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07375__I _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08871_ _02503_ _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07822_ _01291_ _01320_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07753_ _01240_ _01242_ _01287_ _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06704_ _05384_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07684_ _01171_ _01211_ _01212_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09423_ _02319_ _02615_ _02515_ _02309_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06635_ _00083_ _00113_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09354_ _02507_ _02940_ _02937_ _02938_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__08438__A1 _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06566_ _00087_ _00097_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08305_ _01777_ _01886_ _01887_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08989__A2 _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09285_ _02898_ _02900_ _02951_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06497_ _05620_ _05622_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07110__A1 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08236_ _00912_ _00875_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06454__I _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08167_ _01555_ _01631_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07118_ _00559_ _00566_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08098_ _01573_ _01661_ _01587_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07049_ _00432_ _00574_ _00575_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09166__A2 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _03789_ _03790_ _03795_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_76_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06924__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10962_ net101 _04257_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10893_ _04601_ _04696_ _04697_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08844__I _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09626__B1 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09929__A1 _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11376_ _05203_ _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07404__A2 _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10327_ _04053_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05966__A2 _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05708__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10258_ _04006_ _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07168__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10189_ _03935_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08380__A3 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10475__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07340__A1 _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06420_ _05624_ _05627_ _05629_ _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_22_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08754__I _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06351_ _02661_ _05302_ _05126_ _03378_ _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09070_ _02562_ _02717_ _02718_ _02669_ _02675_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_06282_ _05461_ _05493_ _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08840__A1 _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08021_ _01579_ _00211_ _00131_ _01499_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09396__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09972_ _03621_ _03625_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08923_ _02375_ _02250_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08854_ _02477_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07833__I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07805_ _01277_ _01278_ _01329_ _01344_ net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_73_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08785_ _02360_ _02409_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05997_ _01944_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06382__A2 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07736_ _00804_ _00907_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07667_ _00898_ _00131_ _00394_ _01068_ _00891_ _05586_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__A1 _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06618_ _00040_ _00147_ _00148_ _00119_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09406_ _02301_ _02503_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08664__I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07598_ _01075_ _01066_ _01120_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_71_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10218__A1 _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06549_ _00073_ _00080_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09337_ _02858_ _03005_ _03007_ _02928_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10769__A2 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09268_ _02871_ _02870_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_output197_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08219_ _01793_ _01794_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09199_ _02331_ _02385_ _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11230_ net109 net32 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11161_ _04899_ _04988_ _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10112_ net108 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10941__A2 _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06070__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06070__B2 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11092_ _04330_ _04908_ _04913_ _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_103_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10043_ _03689_ _03695_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_76_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07570__A1 _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10945_ _04746_ _04753_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10876_ _04594_ _04628_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07873__A2 _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__A1 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07625__A2 _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11421__A3 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09378__A2 _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11359_ _05144_ _05204_ _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05920_ _03672_ _03727_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08749__I _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05851_ _02976_ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09550__A2 _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10696__A1 _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08570_ _02082_ _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05782_ _02226_ _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07521_ _00840_ _00863_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09302__A2 _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10999__A2 _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07452_ _00944_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06403_ _05556_ _05572_ _05613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07383_ net131 _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09066__A1 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09122_ _02561_ _02598_ _02666_ _02729_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06334_ _05543_ _05485_ _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08813__A1 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09081__A4 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09053_ _02406_ _02407_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06265_ _03444_ _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08004_ _00805_ _00829_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06196_ _05408_ _01987_ _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10254__I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08041__A2 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10923__A2 _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09955_ _03580_ _03582_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08906_ _02377_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08659__I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09886_ _03497_ _03506_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10687__A1 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08837_ _02257_ _02261_ _02417_ _02466_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10687__B2 _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06355__A2 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06179__I _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08768_ _02371_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07719_ _01191_ _01186_ _01201_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_72_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07304__A1 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06107__A2 _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08699_ _02315_ _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10730_ _04437_ _04449_ _04520_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05811__I _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10661_ _04192_ _04446_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09057__A1 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06128__B _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10592_ _04370_ _04371_ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_40_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07607__A2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08280__A2 _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11213_ _05042_ _05044_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10164__I _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11144_ _03861_ _03923_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09780__A2 _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11075_ _03851_ _04231_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput130 b_operand[7] net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10026_ _02292_ _02310_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06346__A2 _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10928_ _04655_ _04736_ net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09048__A1 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10859_ _04580_ _04631_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09048__B2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09599__A2 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06050_ _03063_ _04506_ _05136_ _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11158__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10074__I _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10905__A2 _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07782__A1 _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06952_ _02216_ _02748_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09740_ _02264_ _03351_ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

